module ALU( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [31:0] io_A, // @[:@6.4]
  input  [31:0] io_B, // @[:@6.4]
  input  [3:0]  io_opcode, // @[:@6.4]
  output [31:0] io_out, // @[:@6.4]
  output        io_flagZero // @[:@6.4]
);
  wire [32:0] _T_28; // @[ALU.scala 33:32:@8.4]
  wire [31:0] _T_29; // @[ALU.scala 33:32:@9.4]
  wire [32:0] _T_30; // @[ALU.scala 34:32:@10.4]
  wire [32:0] _T_31; // @[ALU.scala 34:32:@11.4]
  wire [31:0] _T_32; // @[ALU.scala 34:32:@12.4]
  wire [31:0] _T_33; // @[ALU.scala 38:32:@13.4]
  wire [31:0] _T_34; // @[ALU.scala 38:46:@14.4]
  wire  _T_35; // @[ALU.scala 38:39:@15.4]
  wire  _T_36; // @[ALU.scala 39:32:@16.4]
  wire [31:0] _T_37; // @[ALU.scala 40:32:@17.4]
  wire [31:0] _T_38; // @[ALU.scala 41:32:@18.4]
  wire [31:0] _T_39; // @[ALU.scala 42:32:@19.4]
  wire  _T_40; // @[Mux.scala 46:19:@20.4]
  wire [31:0] _T_41; // @[Mux.scala 46:16:@21.4]
  wire  _T_42; // @[Mux.scala 46:19:@22.4]
  wire [31:0] _T_43; // @[Mux.scala 46:16:@23.4]
  wire  _T_44; // @[Mux.scala 46:19:@24.4]
  wire [31:0] _T_45; // @[Mux.scala 46:16:@25.4]
  wire  _T_46; // @[Mux.scala 46:19:@26.4]
  wire [31:0] _T_47; // @[Mux.scala 46:16:@27.4]
  wire  _T_48; // @[Mux.scala 46:19:@28.4]
  wire [31:0] _T_49; // @[Mux.scala 46:16:@29.4]
  wire  _T_50; // @[Mux.scala 46:19:@30.4]
  wire [31:0] _T_51; // @[Mux.scala 46:16:@31.4]
  wire  _T_52; // @[Mux.scala 46:19:@32.4]
  wire [31:0] _T_53; // @[Mux.scala 46:16:@33.4]
  wire  _T_54; // @[Mux.scala 46:19:@34.4]
  assign _T_28 = io_A + io_B; // @[ALU.scala 33:32:@8.4]
  assign _T_29 = io_A + io_B; // @[ALU.scala 33:32:@9.4]
  assign _T_30 = io_A - io_B; // @[ALU.scala 34:32:@10.4]
  assign _T_31 = $unsigned(_T_30); // @[ALU.scala 34:32:@11.4]
  assign _T_32 = _T_31[31:0]; // @[ALU.scala 34:32:@12.4]
  assign _T_33 = $signed(io_A); // @[ALU.scala 38:32:@13.4]
  assign _T_34 = $signed(io_B); // @[ALU.scala 38:46:@14.4]
  assign _T_35 = $signed(_T_33) < $signed(_T_34); // @[ALU.scala 38:39:@15.4]
  assign _T_36 = io_A < io_B; // @[ALU.scala 39:32:@16.4]
  assign _T_37 = io_A & io_B; // @[ALU.scala 40:32:@17.4]
  assign _T_38 = io_A | io_B; // @[ALU.scala 41:32:@18.4]
  assign _T_39 = io_A ^ io_B; // @[ALU.scala 42:32:@19.4]
  assign _T_40 = 4'ha == io_opcode; // @[Mux.scala 46:19:@20.4]
  assign _T_41 = _T_40 ? io_A : io_B; // @[Mux.scala 46:16:@21.4]
  assign _T_42 = 4'h4 == io_opcode; // @[Mux.scala 46:19:@22.4]
  assign _T_43 = _T_42 ? _T_39 : _T_41; // @[Mux.scala 46:16:@23.4]
  assign _T_44 = 4'h3 == io_opcode; // @[Mux.scala 46:19:@24.4]
  assign _T_45 = _T_44 ? _T_38 : _T_43; // @[Mux.scala 46:16:@25.4]
  assign _T_46 = 4'h2 == io_opcode; // @[Mux.scala 46:19:@26.4]
  assign _T_47 = _T_46 ? _T_37 : _T_45; // @[Mux.scala 46:16:@27.4]
  assign _T_48 = 4'h7 == io_opcode; // @[Mux.scala 46:19:@28.4]
  assign _T_49 = _T_48 ? {{31'd0}, _T_36} : _T_47; // @[Mux.scala 46:16:@29.4]
  assign _T_50 = 4'h5 == io_opcode; // @[Mux.scala 46:19:@30.4]
  assign _T_51 = _T_50 ? {{31'd0}, _T_35} : _T_49; // @[Mux.scala 46:16:@31.4]
  assign _T_52 = 4'h1 == io_opcode; // @[Mux.scala 46:19:@32.4]
  assign _T_53 = _T_52 ? _T_32 : _T_51; // @[Mux.scala 46:16:@33.4]
  assign _T_54 = 4'h0 == io_opcode; // @[Mux.scala 46:19:@34.4]
  assign io_out = _T_54 ? _T_29 : _T_53; // @[ALU.scala 32:12:@36.4]
  assign io_flagZero = io_out == 32'h0; // @[ALU.scala 45:17:@38.4]
endmodule
