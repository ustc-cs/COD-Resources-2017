module ALU( // @[:@3.2]
  input  [31:0] io_A, // @[:@6.4]
  input  [31:0] io_B, // @[:@6.4]
  input  [3:0]  io_opcode, // @[:@6.4]
  output [31:0] io_out, // @[:@6.4]
  output        io_flagZero // @[:@6.4]
);
  wire [32:0] _T_29; // @[ALU.scala 34:32:@8.4]
  wire [31:0] _T_30; // @[ALU.scala 34:32:@9.4]
  wire [32:0] _T_31; // @[ALU.scala 35:32:@10.4]
  wire [32:0] _T_32; // @[ALU.scala 35:32:@11.4]
  wire [31:0] _T_33; // @[ALU.scala 35:32:@12.4]
  wire [31:0] _T_34; // @[ALU.scala 39:32:@13.4]
  wire [31:0] _T_35; // @[ALU.scala 39:46:@14.4]
  wire  _T_36; // @[ALU.scala 39:39:@15.4]
  wire  _T_37; // @[ALU.scala 40:32:@16.4]
  wire [31:0] _T_38; // @[ALU.scala 41:32:@17.4]
  wire [31:0] _T_39; // @[ALU.scala 42:32:@18.4]
  wire [31:0] _T_40; // @[ALU.scala 43:32:@19.4]
  wire [31:0] _T_42; // @[ALU.scala 44:26:@21.4]
  wire  _T_43; // @[Mux.scala 46:19:@22.4]
  wire [31:0] _T_44; // @[Mux.scala 46:16:@23.4]
  wire  _T_45; // @[Mux.scala 46:19:@24.4]
  wire [31:0] _T_46; // @[Mux.scala 46:16:@25.4]
  wire  _T_47; // @[Mux.scala 46:19:@26.4]
  wire [31:0] _T_48; // @[Mux.scala 46:16:@27.4]
  wire  _T_49; // @[Mux.scala 46:19:@28.4]
  wire [31:0] _T_50; // @[Mux.scala 46:16:@29.4]
  wire  _T_51; // @[Mux.scala 46:19:@30.4]
  wire [31:0] _T_52; // @[Mux.scala 46:16:@31.4]
  wire  _T_53; // @[Mux.scala 46:19:@32.4]
  wire [31:0] _T_54; // @[Mux.scala 46:16:@33.4]
  wire  _T_55; // @[Mux.scala 46:19:@34.4]
  wire [31:0] _T_56; // @[Mux.scala 46:16:@35.4]
  wire  _T_57; // @[Mux.scala 46:19:@36.4]
  wire [31:0] _T_58; // @[Mux.scala 46:16:@37.4]
  wire  _T_59; // @[Mux.scala 46:19:@38.4]
  assign _T_29 = io_A + io_B; // @[ALU.scala 34:32:@8.4]
  assign _T_30 = io_A + io_B; // @[ALU.scala 34:32:@9.4]
  assign _T_31 = io_A - io_B; // @[ALU.scala 35:32:@10.4]
  assign _T_32 = $unsigned(_T_31); // @[ALU.scala 35:32:@11.4]
  assign _T_33 = _T_32[31:0]; // @[ALU.scala 35:32:@12.4]
  assign _T_34 = $signed(io_A); // @[ALU.scala 39:32:@13.4]
  assign _T_35 = $signed(io_B); // @[ALU.scala 39:46:@14.4]
  assign _T_36 = $signed(_T_34) < $signed(_T_35); // @[ALU.scala 39:39:@15.4]
  assign _T_37 = io_A < io_B; // @[ALU.scala 40:32:@16.4]
  assign _T_38 = io_A & io_B; // @[ALU.scala 41:32:@17.4]
  assign _T_39 = io_A | io_B; // @[ALU.scala 42:32:@18.4]
  assign _T_40 = io_A ^ io_B; // @[ALU.scala 43:32:@19.4]
  assign _T_42 = ~ _T_40; // @[ALU.scala 44:26:@21.4]
  assign _T_43 = 4'ha == io_opcode; // @[Mux.scala 46:19:@22.4]
  assign _T_44 = _T_43 ? io_A : io_B; // @[Mux.scala 46:16:@23.4]
  assign _T_45 = 4'hc == io_opcode; // @[Mux.scala 46:19:@24.4]
  assign _T_46 = _T_45 ? _T_42 : _T_44; // @[Mux.scala 46:16:@25.4]
  assign _T_47 = 4'h4 == io_opcode; // @[Mux.scala 46:19:@26.4]
  assign _T_48 = _T_47 ? _T_40 : _T_46; // @[Mux.scala 46:16:@27.4]
  assign _T_49 = 4'h3 == io_opcode; // @[Mux.scala 46:19:@28.4]
  assign _T_50 = _T_49 ? _T_39 : _T_48; // @[Mux.scala 46:16:@29.4]
  assign _T_51 = 4'h2 == io_opcode; // @[Mux.scala 46:19:@30.4]
  assign _T_52 = _T_51 ? _T_38 : _T_50; // @[Mux.scala 46:16:@31.4]
  assign _T_53 = 4'h7 == io_opcode; // @[Mux.scala 46:19:@32.4]
  assign _T_54 = _T_53 ? {{31'd0}, _T_37} : _T_52; // @[Mux.scala 46:16:@33.4]
  assign _T_55 = 4'h5 == io_opcode; // @[Mux.scala 46:19:@34.4]
  assign _T_56 = _T_55 ? {{31'd0}, _T_36} : _T_54; // @[Mux.scala 46:16:@35.4]
  assign _T_57 = 4'h1 == io_opcode; // @[Mux.scala 46:19:@36.4]
  assign _T_58 = _T_57 ? _T_33 : _T_56; // @[Mux.scala 46:16:@37.4]
  assign _T_59 = 4'h0 == io_opcode; // @[Mux.scala 46:19:@38.4]
  assign io_out = _T_59 ? _T_30 : _T_58; // @[ALU.scala 33:12:@40.4]
  assign io_flagZero = io_out == 32'h0; // @[ALU.scala 47:17:@42.4]
endmodule
module RegFile( // @[:@44.2]
  input         clock, // @[:@45.4]
  input         reset, // @[:@46.4]
  input  [4:0]  io_ra_a, // @[:@47.4]
  input  [4:0]  io_ra_b, // @[:@47.4]
  input  [4:0]  io_wa, // @[:@47.4]
  input  [31:0] io_wd, // @[:@47.4]
  output [31:0] io_rd_a, // @[:@47.4]
  output [31:0] io_rd_b, // @[:@47.4]
  input         io_RegWrite, // @[:@47.4]
  input  [4:0]  io_ra_c, // @[:@47.4]
  output [31:0] io_rd_c // @[:@47.4]
);
  reg [31:0] regs_0; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_0;
  reg [31:0] regs_1; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_1;
  reg [31:0] regs_2; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_2;
  reg [31:0] regs_3; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_3;
  reg [31:0] regs_4; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_4;
  reg [31:0] regs_5; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_5;
  reg [31:0] regs_6; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_6;
  reg [31:0] regs_7; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_7;
  reg [31:0] regs_8; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_8;
  reg [31:0] regs_9; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_9;
  reg [31:0] regs_10; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_10;
  reg [31:0] regs_11; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_11;
  reg [31:0] regs_12; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_12;
  reg [31:0] regs_13; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_13;
  reg [31:0] regs_14; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_14;
  reg [31:0] regs_15; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_15;
  reg [31:0] regs_16; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_16;
  reg [31:0] regs_17; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_17;
  reg [31:0] regs_18; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_18;
  reg [31:0] regs_19; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_19;
  reg [31:0] regs_20; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_20;
  reg [31:0] regs_21; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_21;
  reg [31:0] regs_22; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_22;
  reg [31:0] regs_23; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_23;
  reg [31:0] regs_24; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_24;
  reg [31:0] regs_25; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_25;
  reg [31:0] regs_26; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_26;
  reg [31:0] regs_27; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_27;
  reg [31:0] regs_28; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_28;
  reg [31:0] regs_29; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_29;
  reg [31:0] regs_30; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_30;
  reg [31:0] regs_31; // @[RegFile.scala 21:23:@82.4]
  reg [31:0] _RAND_31;
  wire  _T_262; // @[RegFile.scala 23:21:@83.4]
  wire  _T_263; // @[RegFile.scala 23:34:@84.4]
  wire [31:0] _GEN_0; // @[RegFile.scala 23:50:@85.4]
  wire  _T_265; // @[RegFile.scala 23:21:@88.4]
  wire  _T_266; // @[RegFile.scala 23:34:@89.4]
  wire [31:0] _GEN_1; // @[RegFile.scala 23:50:@90.4]
  wire  _T_268; // @[RegFile.scala 23:21:@93.4]
  wire  _T_269; // @[RegFile.scala 23:34:@94.4]
  wire [31:0] _GEN_2; // @[RegFile.scala 23:50:@95.4]
  wire  _T_271; // @[RegFile.scala 23:21:@98.4]
  wire  _T_272; // @[RegFile.scala 23:34:@99.4]
  wire [31:0] _GEN_3; // @[RegFile.scala 23:50:@100.4]
  wire  _T_274; // @[RegFile.scala 23:21:@103.4]
  wire  _T_275; // @[RegFile.scala 23:34:@104.4]
  wire [31:0] _GEN_4; // @[RegFile.scala 23:50:@105.4]
  wire  _T_277; // @[RegFile.scala 23:21:@108.4]
  wire  _T_278; // @[RegFile.scala 23:34:@109.4]
  wire [31:0] _GEN_5; // @[RegFile.scala 23:50:@110.4]
  wire  _T_280; // @[RegFile.scala 23:21:@113.4]
  wire  _T_281; // @[RegFile.scala 23:34:@114.4]
  wire [31:0] _GEN_6; // @[RegFile.scala 23:50:@115.4]
  wire  _T_283; // @[RegFile.scala 23:21:@118.4]
  wire  _T_284; // @[RegFile.scala 23:34:@119.4]
  wire [31:0] _GEN_7; // @[RegFile.scala 23:50:@120.4]
  wire  _T_286; // @[RegFile.scala 23:21:@123.4]
  wire  _T_287; // @[RegFile.scala 23:34:@124.4]
  wire [31:0] _GEN_8; // @[RegFile.scala 23:50:@125.4]
  wire  _T_289; // @[RegFile.scala 23:21:@128.4]
  wire  _T_290; // @[RegFile.scala 23:34:@129.4]
  wire [31:0] _GEN_9; // @[RegFile.scala 23:50:@130.4]
  wire  _T_292; // @[RegFile.scala 23:21:@133.4]
  wire  _T_293; // @[RegFile.scala 23:34:@134.4]
  wire [31:0] _GEN_10; // @[RegFile.scala 23:50:@135.4]
  wire  _T_295; // @[RegFile.scala 23:21:@138.4]
  wire  _T_296; // @[RegFile.scala 23:34:@139.4]
  wire [31:0] _GEN_11; // @[RegFile.scala 23:50:@140.4]
  wire  _T_298; // @[RegFile.scala 23:21:@143.4]
  wire  _T_299; // @[RegFile.scala 23:34:@144.4]
  wire [31:0] _GEN_12; // @[RegFile.scala 23:50:@145.4]
  wire  _T_301; // @[RegFile.scala 23:21:@148.4]
  wire  _T_302; // @[RegFile.scala 23:34:@149.4]
  wire [31:0] _GEN_13; // @[RegFile.scala 23:50:@150.4]
  wire  _T_304; // @[RegFile.scala 23:21:@153.4]
  wire  _T_305; // @[RegFile.scala 23:34:@154.4]
  wire [31:0] _GEN_14; // @[RegFile.scala 23:50:@155.4]
  wire  _T_307; // @[RegFile.scala 23:21:@158.4]
  wire  _T_308; // @[RegFile.scala 23:34:@159.4]
  wire [31:0] _GEN_15; // @[RegFile.scala 23:50:@160.4]
  wire  _T_310; // @[RegFile.scala 23:21:@163.4]
  wire  _T_311; // @[RegFile.scala 23:34:@164.4]
  wire [31:0] _GEN_16; // @[RegFile.scala 23:50:@165.4]
  wire  _T_313; // @[RegFile.scala 23:21:@168.4]
  wire  _T_314; // @[RegFile.scala 23:34:@169.4]
  wire [31:0] _GEN_17; // @[RegFile.scala 23:50:@170.4]
  wire  _T_316; // @[RegFile.scala 23:21:@173.4]
  wire  _T_317; // @[RegFile.scala 23:34:@174.4]
  wire [31:0] _GEN_18; // @[RegFile.scala 23:50:@175.4]
  wire  _T_319; // @[RegFile.scala 23:21:@178.4]
  wire  _T_320; // @[RegFile.scala 23:34:@179.4]
  wire [31:0] _GEN_19; // @[RegFile.scala 23:50:@180.4]
  wire  _T_322; // @[RegFile.scala 23:21:@183.4]
  wire  _T_323; // @[RegFile.scala 23:34:@184.4]
  wire [31:0] _GEN_20; // @[RegFile.scala 23:50:@185.4]
  wire  _T_325; // @[RegFile.scala 23:21:@188.4]
  wire  _T_326; // @[RegFile.scala 23:34:@189.4]
  wire [31:0] _GEN_21; // @[RegFile.scala 23:50:@190.4]
  wire  _T_328; // @[RegFile.scala 23:21:@193.4]
  wire  _T_329; // @[RegFile.scala 23:34:@194.4]
  wire [31:0] _GEN_22; // @[RegFile.scala 23:50:@195.4]
  wire  _T_331; // @[RegFile.scala 23:21:@198.4]
  wire  _T_332; // @[RegFile.scala 23:34:@199.4]
  wire [31:0] _GEN_23; // @[RegFile.scala 23:50:@200.4]
  wire  _T_334; // @[RegFile.scala 23:21:@203.4]
  wire  _T_335; // @[RegFile.scala 23:34:@204.4]
  wire [31:0] _GEN_24; // @[RegFile.scala 23:50:@205.4]
  wire  _T_337; // @[RegFile.scala 23:21:@208.4]
  wire  _T_338; // @[RegFile.scala 23:34:@209.4]
  wire [31:0] _GEN_25; // @[RegFile.scala 23:50:@210.4]
  wire  _T_340; // @[RegFile.scala 23:21:@213.4]
  wire  _T_341; // @[RegFile.scala 23:34:@214.4]
  wire [31:0] _GEN_26; // @[RegFile.scala 23:50:@215.4]
  wire  _T_343; // @[RegFile.scala 23:21:@218.4]
  wire  _T_344; // @[RegFile.scala 23:34:@219.4]
  wire [31:0] _GEN_27; // @[RegFile.scala 23:50:@220.4]
  wire  _T_346; // @[RegFile.scala 23:21:@223.4]
  wire  _T_347; // @[RegFile.scala 23:34:@224.4]
  wire [31:0] _GEN_28; // @[RegFile.scala 23:50:@225.4]
  wire  _T_349; // @[RegFile.scala 23:21:@228.4]
  wire  _T_350; // @[RegFile.scala 23:34:@229.4]
  wire [31:0] _GEN_29; // @[RegFile.scala 23:50:@230.4]
  wire  _T_352; // @[RegFile.scala 23:21:@233.4]
  wire  _T_353; // @[RegFile.scala 23:34:@234.4]
  wire [31:0] _GEN_30; // @[RegFile.scala 23:50:@235.4]
  wire  _T_355; // @[RegFile.scala 23:21:@238.4]
  wire  _T_356; // @[RegFile.scala 23:34:@239.4]
  wire [31:0] _GEN_31; // @[RegFile.scala 23:50:@240.4]
  wire  raZero; // @[RegFile.scala 33:27:@243.4]
  wire  rbZero; // @[RegFile.scala 34:27:@244.4]
  wire  rcZero; // @[RegFile.scala 35:27:@245.4]
  wire [31:0] _GEN_33; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_34; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_35; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_36; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_37; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_38; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_39; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_40; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_41; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_42; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_43; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_44; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_45; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_46; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_47; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_48; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_49; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_50; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_51; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_52; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_53; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_54; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_55; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_56; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_57; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_58; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_59; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_60; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_61; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_62; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_63; // @[RegFile.scala 36:19:@246.4]
  wire [31:0] _GEN_65; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_66; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_67; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_68; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_69; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_70; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_71; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_72; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_73; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_74; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_75; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_76; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_77; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_78; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_79; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_80; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_81; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_82; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_83; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_84; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_85; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_86; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_87; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_88; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_89; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_90; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_91; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_92; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_93; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_94; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_95; // @[RegFile.scala 37:19:@248.4]
  wire [31:0] _GEN_97; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_98; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_99; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_100; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_101; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_102; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_103; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_104; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_105; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_106; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_107; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_108; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_109; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_110; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_111; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_112; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_113; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_114; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_115; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_116; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_117; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_118; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_119; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_120; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_121; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_122; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_123; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_124; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_125; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_126; // @[RegFile.scala 38:19:@250.4]
  wire [31:0] _GEN_127; // @[RegFile.scala 38:19:@250.4]
  assign _T_262 = io_wa == 5'h0; // @[RegFile.scala 23:21:@83.4]
  assign _T_263 = _T_262 & io_RegWrite; // @[RegFile.scala 23:34:@84.4]
  assign _GEN_0 = _T_263 ? io_wd : regs_0; // @[RegFile.scala 23:50:@85.4]
  assign _T_265 = io_wa == 5'h1; // @[RegFile.scala 23:21:@88.4]
  assign _T_266 = _T_265 & io_RegWrite; // @[RegFile.scala 23:34:@89.4]
  assign _GEN_1 = _T_266 ? io_wd : regs_1; // @[RegFile.scala 23:50:@90.4]
  assign _T_268 = io_wa == 5'h2; // @[RegFile.scala 23:21:@93.4]
  assign _T_269 = _T_268 & io_RegWrite; // @[RegFile.scala 23:34:@94.4]
  assign _GEN_2 = _T_269 ? io_wd : regs_2; // @[RegFile.scala 23:50:@95.4]
  assign _T_271 = io_wa == 5'h3; // @[RegFile.scala 23:21:@98.4]
  assign _T_272 = _T_271 & io_RegWrite; // @[RegFile.scala 23:34:@99.4]
  assign _GEN_3 = _T_272 ? io_wd : regs_3; // @[RegFile.scala 23:50:@100.4]
  assign _T_274 = io_wa == 5'h4; // @[RegFile.scala 23:21:@103.4]
  assign _T_275 = _T_274 & io_RegWrite; // @[RegFile.scala 23:34:@104.4]
  assign _GEN_4 = _T_275 ? io_wd : regs_4; // @[RegFile.scala 23:50:@105.4]
  assign _T_277 = io_wa == 5'h5; // @[RegFile.scala 23:21:@108.4]
  assign _T_278 = _T_277 & io_RegWrite; // @[RegFile.scala 23:34:@109.4]
  assign _GEN_5 = _T_278 ? io_wd : regs_5; // @[RegFile.scala 23:50:@110.4]
  assign _T_280 = io_wa == 5'h6; // @[RegFile.scala 23:21:@113.4]
  assign _T_281 = _T_280 & io_RegWrite; // @[RegFile.scala 23:34:@114.4]
  assign _GEN_6 = _T_281 ? io_wd : regs_6; // @[RegFile.scala 23:50:@115.4]
  assign _T_283 = io_wa == 5'h7; // @[RegFile.scala 23:21:@118.4]
  assign _T_284 = _T_283 & io_RegWrite; // @[RegFile.scala 23:34:@119.4]
  assign _GEN_7 = _T_284 ? io_wd : regs_7; // @[RegFile.scala 23:50:@120.4]
  assign _T_286 = io_wa == 5'h8; // @[RegFile.scala 23:21:@123.4]
  assign _T_287 = _T_286 & io_RegWrite; // @[RegFile.scala 23:34:@124.4]
  assign _GEN_8 = _T_287 ? io_wd : regs_8; // @[RegFile.scala 23:50:@125.4]
  assign _T_289 = io_wa == 5'h9; // @[RegFile.scala 23:21:@128.4]
  assign _T_290 = _T_289 & io_RegWrite; // @[RegFile.scala 23:34:@129.4]
  assign _GEN_9 = _T_290 ? io_wd : regs_9; // @[RegFile.scala 23:50:@130.4]
  assign _T_292 = io_wa == 5'ha; // @[RegFile.scala 23:21:@133.4]
  assign _T_293 = _T_292 & io_RegWrite; // @[RegFile.scala 23:34:@134.4]
  assign _GEN_10 = _T_293 ? io_wd : regs_10; // @[RegFile.scala 23:50:@135.4]
  assign _T_295 = io_wa == 5'hb; // @[RegFile.scala 23:21:@138.4]
  assign _T_296 = _T_295 & io_RegWrite; // @[RegFile.scala 23:34:@139.4]
  assign _GEN_11 = _T_296 ? io_wd : regs_11; // @[RegFile.scala 23:50:@140.4]
  assign _T_298 = io_wa == 5'hc; // @[RegFile.scala 23:21:@143.4]
  assign _T_299 = _T_298 & io_RegWrite; // @[RegFile.scala 23:34:@144.4]
  assign _GEN_12 = _T_299 ? io_wd : regs_12; // @[RegFile.scala 23:50:@145.4]
  assign _T_301 = io_wa == 5'hd; // @[RegFile.scala 23:21:@148.4]
  assign _T_302 = _T_301 & io_RegWrite; // @[RegFile.scala 23:34:@149.4]
  assign _GEN_13 = _T_302 ? io_wd : regs_13; // @[RegFile.scala 23:50:@150.4]
  assign _T_304 = io_wa == 5'he; // @[RegFile.scala 23:21:@153.4]
  assign _T_305 = _T_304 & io_RegWrite; // @[RegFile.scala 23:34:@154.4]
  assign _GEN_14 = _T_305 ? io_wd : regs_14; // @[RegFile.scala 23:50:@155.4]
  assign _T_307 = io_wa == 5'hf; // @[RegFile.scala 23:21:@158.4]
  assign _T_308 = _T_307 & io_RegWrite; // @[RegFile.scala 23:34:@159.4]
  assign _GEN_15 = _T_308 ? io_wd : regs_15; // @[RegFile.scala 23:50:@160.4]
  assign _T_310 = io_wa == 5'h10; // @[RegFile.scala 23:21:@163.4]
  assign _T_311 = _T_310 & io_RegWrite; // @[RegFile.scala 23:34:@164.4]
  assign _GEN_16 = _T_311 ? io_wd : regs_16; // @[RegFile.scala 23:50:@165.4]
  assign _T_313 = io_wa == 5'h11; // @[RegFile.scala 23:21:@168.4]
  assign _T_314 = _T_313 & io_RegWrite; // @[RegFile.scala 23:34:@169.4]
  assign _GEN_17 = _T_314 ? io_wd : regs_17; // @[RegFile.scala 23:50:@170.4]
  assign _T_316 = io_wa == 5'h12; // @[RegFile.scala 23:21:@173.4]
  assign _T_317 = _T_316 & io_RegWrite; // @[RegFile.scala 23:34:@174.4]
  assign _GEN_18 = _T_317 ? io_wd : regs_18; // @[RegFile.scala 23:50:@175.4]
  assign _T_319 = io_wa == 5'h13; // @[RegFile.scala 23:21:@178.4]
  assign _T_320 = _T_319 & io_RegWrite; // @[RegFile.scala 23:34:@179.4]
  assign _GEN_19 = _T_320 ? io_wd : regs_19; // @[RegFile.scala 23:50:@180.4]
  assign _T_322 = io_wa == 5'h14; // @[RegFile.scala 23:21:@183.4]
  assign _T_323 = _T_322 & io_RegWrite; // @[RegFile.scala 23:34:@184.4]
  assign _GEN_20 = _T_323 ? io_wd : regs_20; // @[RegFile.scala 23:50:@185.4]
  assign _T_325 = io_wa == 5'h15; // @[RegFile.scala 23:21:@188.4]
  assign _T_326 = _T_325 & io_RegWrite; // @[RegFile.scala 23:34:@189.4]
  assign _GEN_21 = _T_326 ? io_wd : regs_21; // @[RegFile.scala 23:50:@190.4]
  assign _T_328 = io_wa == 5'h16; // @[RegFile.scala 23:21:@193.4]
  assign _T_329 = _T_328 & io_RegWrite; // @[RegFile.scala 23:34:@194.4]
  assign _GEN_22 = _T_329 ? io_wd : regs_22; // @[RegFile.scala 23:50:@195.4]
  assign _T_331 = io_wa == 5'h17; // @[RegFile.scala 23:21:@198.4]
  assign _T_332 = _T_331 & io_RegWrite; // @[RegFile.scala 23:34:@199.4]
  assign _GEN_23 = _T_332 ? io_wd : regs_23; // @[RegFile.scala 23:50:@200.4]
  assign _T_334 = io_wa == 5'h18; // @[RegFile.scala 23:21:@203.4]
  assign _T_335 = _T_334 & io_RegWrite; // @[RegFile.scala 23:34:@204.4]
  assign _GEN_24 = _T_335 ? io_wd : regs_24; // @[RegFile.scala 23:50:@205.4]
  assign _T_337 = io_wa == 5'h19; // @[RegFile.scala 23:21:@208.4]
  assign _T_338 = _T_337 & io_RegWrite; // @[RegFile.scala 23:34:@209.4]
  assign _GEN_25 = _T_338 ? io_wd : regs_25; // @[RegFile.scala 23:50:@210.4]
  assign _T_340 = io_wa == 5'h1a; // @[RegFile.scala 23:21:@213.4]
  assign _T_341 = _T_340 & io_RegWrite; // @[RegFile.scala 23:34:@214.4]
  assign _GEN_26 = _T_341 ? io_wd : regs_26; // @[RegFile.scala 23:50:@215.4]
  assign _T_343 = io_wa == 5'h1b; // @[RegFile.scala 23:21:@218.4]
  assign _T_344 = _T_343 & io_RegWrite; // @[RegFile.scala 23:34:@219.4]
  assign _GEN_27 = _T_344 ? io_wd : regs_27; // @[RegFile.scala 23:50:@220.4]
  assign _T_346 = io_wa == 5'h1c; // @[RegFile.scala 23:21:@223.4]
  assign _T_347 = _T_346 & io_RegWrite; // @[RegFile.scala 23:34:@224.4]
  assign _GEN_28 = _T_347 ? io_wd : regs_28; // @[RegFile.scala 23:50:@225.4]
  assign _T_349 = io_wa == 5'h1d; // @[RegFile.scala 23:21:@228.4]
  assign _T_350 = _T_349 & io_RegWrite; // @[RegFile.scala 23:34:@229.4]
  assign _GEN_29 = _T_350 ? io_wd : regs_29; // @[RegFile.scala 23:50:@230.4]
  assign _T_352 = io_wa == 5'h1e; // @[RegFile.scala 23:21:@233.4]
  assign _T_353 = _T_352 & io_RegWrite; // @[RegFile.scala 23:34:@234.4]
  assign _GEN_30 = _T_353 ? io_wd : regs_30; // @[RegFile.scala 23:50:@235.4]
  assign _T_355 = io_wa == 5'h1f; // @[RegFile.scala 23:21:@238.4]
  assign _T_356 = _T_355 & io_RegWrite; // @[RegFile.scala 23:34:@239.4]
  assign _GEN_31 = _T_356 ? io_wd : regs_31; // @[RegFile.scala 23:50:@240.4]
  assign raZero = io_ra_a == 5'h0; // @[RegFile.scala 33:27:@243.4]
  assign rbZero = io_ra_b == 5'h0; // @[RegFile.scala 34:27:@244.4]
  assign rcZero = io_ra_c == 5'h0; // @[RegFile.scala 35:27:@245.4]
  assign _GEN_33 = 5'h1 == io_ra_a ? regs_1 : regs_0; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_34 = 5'h2 == io_ra_a ? regs_2 : _GEN_33; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_35 = 5'h3 == io_ra_a ? regs_3 : _GEN_34; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_36 = 5'h4 == io_ra_a ? regs_4 : _GEN_35; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_37 = 5'h5 == io_ra_a ? regs_5 : _GEN_36; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_38 = 5'h6 == io_ra_a ? regs_6 : _GEN_37; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_39 = 5'h7 == io_ra_a ? regs_7 : _GEN_38; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_40 = 5'h8 == io_ra_a ? regs_8 : _GEN_39; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_41 = 5'h9 == io_ra_a ? regs_9 : _GEN_40; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_42 = 5'ha == io_ra_a ? regs_10 : _GEN_41; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_43 = 5'hb == io_ra_a ? regs_11 : _GEN_42; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_44 = 5'hc == io_ra_a ? regs_12 : _GEN_43; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_45 = 5'hd == io_ra_a ? regs_13 : _GEN_44; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_46 = 5'he == io_ra_a ? regs_14 : _GEN_45; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_47 = 5'hf == io_ra_a ? regs_15 : _GEN_46; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_48 = 5'h10 == io_ra_a ? regs_16 : _GEN_47; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_49 = 5'h11 == io_ra_a ? regs_17 : _GEN_48; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_50 = 5'h12 == io_ra_a ? regs_18 : _GEN_49; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_51 = 5'h13 == io_ra_a ? regs_19 : _GEN_50; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_52 = 5'h14 == io_ra_a ? regs_20 : _GEN_51; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_53 = 5'h15 == io_ra_a ? regs_21 : _GEN_52; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_54 = 5'h16 == io_ra_a ? regs_22 : _GEN_53; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_55 = 5'h17 == io_ra_a ? regs_23 : _GEN_54; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_56 = 5'h18 == io_ra_a ? regs_24 : _GEN_55; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_57 = 5'h19 == io_ra_a ? regs_25 : _GEN_56; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_58 = 5'h1a == io_ra_a ? regs_26 : _GEN_57; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_59 = 5'h1b == io_ra_a ? regs_27 : _GEN_58; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_60 = 5'h1c == io_ra_a ? regs_28 : _GEN_59; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_61 = 5'h1d == io_ra_a ? regs_29 : _GEN_60; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_62 = 5'h1e == io_ra_a ? regs_30 : _GEN_61; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_63 = 5'h1f == io_ra_a ? regs_31 : _GEN_62; // @[RegFile.scala 36:19:@246.4]
  assign _GEN_65 = 5'h1 == io_ra_b ? regs_1 : regs_0; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_66 = 5'h2 == io_ra_b ? regs_2 : _GEN_65; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_67 = 5'h3 == io_ra_b ? regs_3 : _GEN_66; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_68 = 5'h4 == io_ra_b ? regs_4 : _GEN_67; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_69 = 5'h5 == io_ra_b ? regs_5 : _GEN_68; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_70 = 5'h6 == io_ra_b ? regs_6 : _GEN_69; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_71 = 5'h7 == io_ra_b ? regs_7 : _GEN_70; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_72 = 5'h8 == io_ra_b ? regs_8 : _GEN_71; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_73 = 5'h9 == io_ra_b ? regs_9 : _GEN_72; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_74 = 5'ha == io_ra_b ? regs_10 : _GEN_73; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_75 = 5'hb == io_ra_b ? regs_11 : _GEN_74; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_76 = 5'hc == io_ra_b ? regs_12 : _GEN_75; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_77 = 5'hd == io_ra_b ? regs_13 : _GEN_76; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_78 = 5'he == io_ra_b ? regs_14 : _GEN_77; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_79 = 5'hf == io_ra_b ? regs_15 : _GEN_78; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_80 = 5'h10 == io_ra_b ? regs_16 : _GEN_79; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_81 = 5'h11 == io_ra_b ? regs_17 : _GEN_80; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_82 = 5'h12 == io_ra_b ? regs_18 : _GEN_81; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_83 = 5'h13 == io_ra_b ? regs_19 : _GEN_82; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_84 = 5'h14 == io_ra_b ? regs_20 : _GEN_83; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_85 = 5'h15 == io_ra_b ? regs_21 : _GEN_84; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_86 = 5'h16 == io_ra_b ? regs_22 : _GEN_85; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_87 = 5'h17 == io_ra_b ? regs_23 : _GEN_86; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_88 = 5'h18 == io_ra_b ? regs_24 : _GEN_87; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_89 = 5'h19 == io_ra_b ? regs_25 : _GEN_88; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_90 = 5'h1a == io_ra_b ? regs_26 : _GEN_89; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_91 = 5'h1b == io_ra_b ? regs_27 : _GEN_90; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_92 = 5'h1c == io_ra_b ? regs_28 : _GEN_91; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_93 = 5'h1d == io_ra_b ? regs_29 : _GEN_92; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_94 = 5'h1e == io_ra_b ? regs_30 : _GEN_93; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_95 = 5'h1f == io_ra_b ? regs_31 : _GEN_94; // @[RegFile.scala 37:19:@248.4]
  assign _GEN_97 = 5'h1 == io_ra_c ? regs_1 : regs_0; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_98 = 5'h2 == io_ra_c ? regs_2 : _GEN_97; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_99 = 5'h3 == io_ra_c ? regs_3 : _GEN_98; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_100 = 5'h4 == io_ra_c ? regs_4 : _GEN_99; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_101 = 5'h5 == io_ra_c ? regs_5 : _GEN_100; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_102 = 5'h6 == io_ra_c ? regs_6 : _GEN_101; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_103 = 5'h7 == io_ra_c ? regs_7 : _GEN_102; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_104 = 5'h8 == io_ra_c ? regs_8 : _GEN_103; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_105 = 5'h9 == io_ra_c ? regs_9 : _GEN_104; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_106 = 5'ha == io_ra_c ? regs_10 : _GEN_105; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_107 = 5'hb == io_ra_c ? regs_11 : _GEN_106; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_108 = 5'hc == io_ra_c ? regs_12 : _GEN_107; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_109 = 5'hd == io_ra_c ? regs_13 : _GEN_108; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_110 = 5'he == io_ra_c ? regs_14 : _GEN_109; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_111 = 5'hf == io_ra_c ? regs_15 : _GEN_110; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_112 = 5'h10 == io_ra_c ? regs_16 : _GEN_111; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_113 = 5'h11 == io_ra_c ? regs_17 : _GEN_112; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_114 = 5'h12 == io_ra_c ? regs_18 : _GEN_113; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_115 = 5'h13 == io_ra_c ? regs_19 : _GEN_114; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_116 = 5'h14 == io_ra_c ? regs_20 : _GEN_115; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_117 = 5'h15 == io_ra_c ? regs_21 : _GEN_116; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_118 = 5'h16 == io_ra_c ? regs_22 : _GEN_117; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_119 = 5'h17 == io_ra_c ? regs_23 : _GEN_118; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_120 = 5'h18 == io_ra_c ? regs_24 : _GEN_119; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_121 = 5'h19 == io_ra_c ? regs_25 : _GEN_120; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_122 = 5'h1a == io_ra_c ? regs_26 : _GEN_121; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_123 = 5'h1b == io_ra_c ? regs_27 : _GEN_122; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_124 = 5'h1c == io_ra_c ? regs_28 : _GEN_123; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_125 = 5'h1d == io_ra_c ? regs_29 : _GEN_124; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_126 = 5'h1e == io_ra_c ? regs_30 : _GEN_125; // @[RegFile.scala 38:19:@250.4]
  assign _GEN_127 = 5'h1f == io_ra_c ? regs_31 : _GEN_126; // @[RegFile.scala 38:19:@250.4]
  assign io_rd_a = raZero ? 32'h0 : _GEN_63; // @[RegFile.scala 36:13:@247.4]
  assign io_rd_b = rbZero ? 32'h0 : _GEN_95; // @[RegFile.scala 37:13:@249.4]
  assign io_rd_c = rcZero ? 32'h0 : _GEN_127; // @[RegFile.scala 38:13:@251.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 32'h0;
    end else begin
      if (_T_263) begin
        regs_0 <= io_wd;
      end
    end
    if (reset) begin
      regs_1 <= 32'h0;
    end else begin
      if (_T_266) begin
        regs_1 <= io_wd;
      end
    end
    if (reset) begin
      regs_2 <= 32'h0;
    end else begin
      if (_T_269) begin
        regs_2 <= io_wd;
      end
    end
    if (reset) begin
      regs_3 <= 32'h0;
    end else begin
      if (_T_272) begin
        regs_3 <= io_wd;
      end
    end
    if (reset) begin
      regs_4 <= 32'h0;
    end else begin
      if (_T_275) begin
        regs_4 <= io_wd;
      end
    end
    if (reset) begin
      regs_5 <= 32'h0;
    end else begin
      if (_T_278) begin
        regs_5 <= io_wd;
      end
    end
    if (reset) begin
      regs_6 <= 32'h0;
    end else begin
      if (_T_281) begin
        regs_6 <= io_wd;
      end
    end
    if (reset) begin
      regs_7 <= 32'h0;
    end else begin
      if (_T_284) begin
        regs_7 <= io_wd;
      end
    end
    if (reset) begin
      regs_8 <= 32'h0;
    end else begin
      if (_T_287) begin
        regs_8 <= io_wd;
      end
    end
    if (reset) begin
      regs_9 <= 32'h0;
    end else begin
      if (_T_290) begin
        regs_9 <= io_wd;
      end
    end
    if (reset) begin
      regs_10 <= 32'h0;
    end else begin
      if (_T_293) begin
        regs_10 <= io_wd;
      end
    end
    if (reset) begin
      regs_11 <= 32'h0;
    end else begin
      if (_T_296) begin
        regs_11 <= io_wd;
      end
    end
    if (reset) begin
      regs_12 <= 32'h0;
    end else begin
      if (_T_299) begin
        regs_12 <= io_wd;
      end
    end
    if (reset) begin
      regs_13 <= 32'h0;
    end else begin
      if (_T_302) begin
        regs_13 <= io_wd;
      end
    end
    if (reset) begin
      regs_14 <= 32'h0;
    end else begin
      if (_T_305) begin
        regs_14 <= io_wd;
      end
    end
    if (reset) begin
      regs_15 <= 32'h0;
    end else begin
      if (_T_308) begin
        regs_15 <= io_wd;
      end
    end
    if (reset) begin
      regs_16 <= 32'h0;
    end else begin
      if (_T_311) begin
        regs_16 <= io_wd;
      end
    end
    if (reset) begin
      regs_17 <= 32'h0;
    end else begin
      if (_T_314) begin
        regs_17 <= io_wd;
      end
    end
    if (reset) begin
      regs_18 <= 32'h0;
    end else begin
      if (_T_317) begin
        regs_18 <= io_wd;
      end
    end
    if (reset) begin
      regs_19 <= 32'h0;
    end else begin
      if (_T_320) begin
        regs_19 <= io_wd;
      end
    end
    if (reset) begin
      regs_20 <= 32'h0;
    end else begin
      if (_T_323) begin
        regs_20 <= io_wd;
      end
    end
    if (reset) begin
      regs_21 <= 32'h0;
    end else begin
      if (_T_326) begin
        regs_21 <= io_wd;
      end
    end
    if (reset) begin
      regs_22 <= 32'h0;
    end else begin
      if (_T_329) begin
        regs_22 <= io_wd;
      end
    end
    if (reset) begin
      regs_23 <= 32'h0;
    end else begin
      if (_T_332) begin
        regs_23 <= io_wd;
      end
    end
    if (reset) begin
      regs_24 <= 32'h0;
    end else begin
      if (_T_335) begin
        regs_24 <= io_wd;
      end
    end
    if (reset) begin
      regs_25 <= 32'h0;
    end else begin
      if (_T_338) begin
        regs_25 <= io_wd;
      end
    end
    if (reset) begin
      regs_26 <= 32'h0;
    end else begin
      if (_T_341) begin
        regs_26 <= io_wd;
      end
    end
    if (reset) begin
      regs_27 <= 32'h0;
    end else begin
      if (_T_344) begin
        regs_27 <= io_wd;
      end
    end
    if (reset) begin
      regs_28 <= 32'h0;
    end else begin
      if (_T_347) begin
        regs_28 <= io_wd;
      end
    end
    if (reset) begin
      regs_29 <= 32'h0;
    end else begin
      if (_T_350) begin
        regs_29 <= io_wd;
      end
    end
    if (reset) begin
      regs_30 <= 32'h0;
    end else begin
      if (_T_353) begin
        regs_30 <= io_wd;
      end
    end
    if (reset) begin
      regs_31 <= 32'h0;
    end else begin
      if (_T_356) begin
        regs_31 <= io_wd;
      end
    end
  end
endmodule
module Datapath( // @[:@253.2]
  input         clock, // @[:@254.4]
  input         reset, // @[:@255.4]
  output [31:0] io_ctrl_Inst, // @[:@256.4]
  input         io_ctrl_IRWrite, // @[:@256.4]
  input         io_ctrl_RegDst, // @[:@256.4]
  input         io_ctrl_RegWrite, // @[:@256.4]
  input         io_ctrl_ALUSrcA, // @[:@256.4]
  input  [2:0]  io_ctrl_ALUSrcB, // @[:@256.4]
  input  [3:0]  io_ctrl_ALUOp, // @[:@256.4]
  input  [1:0]  io_ctrl_PCSource, // @[:@256.4]
  input         io_ctrl_PCWriteBEQ, // @[:@256.4]
  input         io_ctrl_PCWriteBNE, // @[:@256.4]
  input         io_ctrl_PCWrite, // @[:@256.4]
  input         io_ctrl_IorD, // @[:@256.4]
  input         io_ctrl_MemWrite, // @[:@256.4]
  input         io_ctrl_MemtoReg, // @[:@256.4]
  input  [31:0] io_mem_mem_rdata, // @[:@256.4]
  output [31:0] io_mem_mem_addr, // @[:@256.4]
  output [31:0] io_mem_mem_wdata, // @[:@256.4]
  output        io_mem_mem_wen, // @[:@256.4]
  output [31:0] io_debug_ir, // @[:@256.4]
  output [31:0] io_debug_mdr, // @[:@256.4]
  output [31:0] io_debug_aluout, // @[:@256.4]
  output [31:0] io_debug_pc, // @[:@256.4]
  input  [4:0]  io_debug_ra_c, // @[:@256.4]
  output [31:0] io_debug_rd_c // @[:@256.4]
);
  wire [31:0] alu_io_A; // @[Datapath.scala 23:21:@258.4]
  wire [31:0] alu_io_B; // @[Datapath.scala 23:21:@258.4]
  wire [3:0] alu_io_opcode; // @[Datapath.scala 23:21:@258.4]
  wire [31:0] alu_io_out; // @[Datapath.scala 23:21:@258.4]
  wire  alu_io_flagZero; // @[Datapath.scala 23:21:@258.4]
  wire  regFile_clock; // @[Datapath.scala 24:25:@261.4]
  wire  regFile_reset; // @[Datapath.scala 24:25:@261.4]
  wire [4:0] regFile_io_ra_a; // @[Datapath.scala 24:25:@261.4]
  wire [4:0] regFile_io_ra_b; // @[Datapath.scala 24:25:@261.4]
  wire [4:0] regFile_io_wa; // @[Datapath.scala 24:25:@261.4]
  wire [31:0] regFile_io_wd; // @[Datapath.scala 24:25:@261.4]
  wire [31:0] regFile_io_rd_a; // @[Datapath.scala 24:25:@261.4]
  wire [31:0] regFile_io_rd_b; // @[Datapath.scala 24:25:@261.4]
  wire  regFile_io_RegWrite; // @[Datapath.scala 24:25:@261.4]
  wire [4:0] regFile_io_ra_c; // @[Datapath.scala 24:25:@261.4]
  wire [31:0] regFile_io_rd_c; // @[Datapath.scala 24:25:@261.4]
  reg [31:0] ir; // @[Datapath.scala 29:21:@264.4]
  reg [31:0] _RAND_0;
  wire [31:0] _GEN_0; // @[Datapath.scala 30:28:@265.4]
  reg [31:0] mdr; // @[Datapath.scala 36:22:@269.4]
  reg [31:0] _RAND_1;
  reg [31:0] aluout; // @[Datapath.scala 39:25:@271.4]
  reg [31:0] _RAND_2;
  reg [31:0] pc; // @[Datapath.scala 42:21:@273.4]
  reg [31:0] _RAND_3;
  wire  _T_77; // @[Datapath.scala 43:32:@274.4]
  wire  _T_79; // @[Datapath.scala 44:36:@275.4]
  wire  _T_80; // @[Datapath.scala 44:32:@276.4]
  wire  _T_81; // @[Datapath.scala 43:55:@277.4]
  wire  _T_82; // @[Datapath.scala 44:55:@278.4]
  wire [3:0] _T_87; // @[Datapath.scala 49:39:@280.6]
  wire [25:0] _T_88; // @[Datapath.scala 49:51:@281.6]
  wire [27:0] _GEN_2; // @[Datapath.scala 49:58:@282.6]
  wire [27:0] _T_89; // @[Datapath.scala 49:58:@282.6]
  wire [31:0] _T_90; // @[Cat.scala 30:58:@283.6]
  wire  _T_91; // @[Mux.scala 46:19:@284.6]
  wire [31:0] _T_92; // @[Mux.scala 46:16:@285.6]
  wire  _T_93; // @[Mux.scala 46:19:@286.6]
  wire [31:0] _T_94; // @[Mux.scala 46:16:@287.6]
  wire  _T_95; // @[Mux.scala 46:19:@288.6]
  wire [31:0] _T_96; // @[Mux.scala 46:16:@289.6]
  wire [31:0] _GEN_1; // @[Datapath.scala 45:31:@279.4]
  wire [4:0] _T_98; // @[Datapath.scala 55:26:@294.4]
  wire [4:0] _T_99; // @[Datapath.scala 56:46:@296.4]
  wire [15:0] _T_111; // @[Datapath.scala 67:32:@305.4]
  wire [15:0] _T_112; // @[Datapath.scala 67:39:@306.4]
  wire [15:0] _T_113; // @[Datapath.scala 67:46:@307.4]
  wire [17:0] _GEN_3; // @[Datapath.scala 68:47:@310.4]
  wire [17:0] _T_116; // @[Datapath.scala 68:47:@310.4]
  wire [17:0] _T_117; // @[Datapath.scala 68:53:@311.4]
  wire [3:0] _GEN_4; // @[Mux.scala 46:19:@313.4]
  wire  _T_119; // @[Mux.scala 46:19:@313.4]
  wire [15:0] _T_120; // @[Mux.scala 46:16:@314.4]
  wire  _T_121; // @[Mux.scala 46:19:@315.4]
  wire [17:0] _T_122; // @[Mux.scala 46:16:@316.4]
  wire  _T_123; // @[Mux.scala 46:19:@317.4]
  wire [17:0] _T_124; // @[Mux.scala 46:16:@318.4]
  wire  _T_125; // @[Mux.scala 46:19:@319.4]
  wire [31:0] _T_126; // @[Mux.scala 46:16:@320.4]
  wire  _T_127; // @[Mux.scala 46:19:@321.4]
  ALU alu ( // @[Datapath.scala 23:21:@258.4]
    .io_A(alu_io_A),
    .io_B(alu_io_B),
    .io_opcode(alu_io_opcode),
    .io_out(alu_io_out),
    .io_flagZero(alu_io_flagZero)
  );
  RegFile regFile ( // @[Datapath.scala 24:25:@261.4]
    .clock(regFile_clock),
    .reset(regFile_reset),
    .io_ra_a(regFile_io_ra_a),
    .io_ra_b(regFile_io_ra_b),
    .io_wa(regFile_io_wa),
    .io_wd(regFile_io_wd),
    .io_rd_a(regFile_io_rd_a),
    .io_rd_b(regFile_io_rd_b),
    .io_RegWrite(regFile_io_RegWrite),
    .io_ra_c(regFile_io_ra_c),
    .io_rd_c(regFile_io_rd_c)
  );
  assign _GEN_0 = io_ctrl_IRWrite ? io_mem_mem_rdata : ir; // @[Datapath.scala 30:28:@265.4]
  assign _T_77 = io_ctrl_PCWriteBEQ & alu_io_flagZero; // @[Datapath.scala 43:32:@274.4]
  assign _T_79 = alu_io_flagZero == 1'h0; // @[Datapath.scala 44:36:@275.4]
  assign _T_80 = io_ctrl_PCWriteBNE & _T_79; // @[Datapath.scala 44:32:@276.4]
  assign _T_81 = _T_77 | _T_80; // @[Datapath.scala 43:55:@277.4]
  assign _T_82 = _T_81 | io_ctrl_PCWrite; // @[Datapath.scala 44:55:@278.4]
  assign _T_87 = pc[31:28]; // @[Datapath.scala 49:39:@280.6]
  assign _T_88 = ir[25:0]; // @[Datapath.scala 49:51:@281.6]
  assign _GEN_2 = {{2'd0}, _T_88}; // @[Datapath.scala 49:58:@282.6]
  assign _T_89 = _GEN_2 << 2; // @[Datapath.scala 49:58:@282.6]
  assign _T_90 = {_T_87,_T_89}; // @[Cat.scala 30:58:@283.6]
  assign _T_91 = 2'h2 == io_ctrl_PCSource; // @[Mux.scala 46:19:@284.6]
  assign _T_92 = _T_91 ? _T_90 : 32'h0; // @[Mux.scala 46:16:@285.6]
  assign _T_93 = 2'h1 == io_ctrl_PCSource; // @[Mux.scala 46:19:@286.6]
  assign _T_94 = _T_93 ? aluout : _T_92; // @[Mux.scala 46:16:@287.6]
  assign _T_95 = 2'h0 == io_ctrl_PCSource; // @[Mux.scala 46:19:@288.6]
  assign _T_96 = _T_95 ? alu_io_out : _T_94; // @[Mux.scala 46:16:@289.6]
  assign _GEN_1 = _T_82 ? _T_96 : pc; // @[Datapath.scala 45:31:@279.4]
  assign _T_98 = ir[20:16]; // @[Datapath.scala 55:26:@294.4]
  assign _T_99 = ir[15:11]; // @[Datapath.scala 56:46:@296.4]
  assign _T_111 = ir[15:0]; // @[Datapath.scala 67:32:@305.4]
  assign _T_112 = $signed(_T_111); // @[Datapath.scala 67:39:@306.4]
  assign _T_113 = $unsigned(_T_112); // @[Datapath.scala 67:46:@307.4]
  assign _GEN_3 = {{2{_T_112[15]}},_T_112}; // @[Datapath.scala 68:47:@310.4]
  assign _T_116 = $signed(_GEN_3) << 2; // @[Datapath.scala 68:47:@310.4]
  assign _T_117 = $unsigned(_T_116); // @[Datapath.scala 68:53:@311.4]
  assign _GEN_4 = {{1'd0}, io_ctrl_ALUSrcB}; // @[Mux.scala 46:19:@313.4]
  assign _T_119 = 4'h4 == _GEN_4; // @[Mux.scala 46:19:@313.4]
  assign _T_120 = _T_119 ? _T_111 : 16'h0; // @[Mux.scala 46:16:@314.4]
  assign _T_121 = 3'h3 == io_ctrl_ALUSrcB; // @[Mux.scala 46:19:@315.4]
  assign _T_122 = _T_121 ? _T_117 : {{2'd0}, _T_120}; // @[Mux.scala 46:16:@316.4]
  assign _T_123 = 3'h2 == io_ctrl_ALUSrcB; // @[Mux.scala 46:19:@317.4]
  assign _T_124 = _T_123 ? {{2'd0}, _T_113} : _T_122; // @[Mux.scala 46:16:@318.4]
  assign _T_125 = 3'h1 == io_ctrl_ALUSrcB; // @[Mux.scala 46:19:@319.4]
  assign _T_126 = _T_125 ? 32'h4 : {{14'd0}, _T_124}; // @[Mux.scala 46:16:@320.4]
  assign _T_127 = 3'h0 == io_ctrl_ALUSrcB; // @[Mux.scala 46:19:@321.4]
  assign io_ctrl_Inst = ir; // @[Datapath.scala 33:18:@268.4]
  assign io_mem_mem_addr = io_ctrl_IorD ? aluout : pc; // @[Datapath.scala 76:22:@326.4]
  assign io_mem_mem_wdata = regFile_io_rd_b; // @[Datapath.scala 77:22:@327.4]
  assign io_mem_mem_wen = io_ctrl_MemWrite; // @[Datapath.scala 78:22:@328.4]
  assign io_debug_ir = ir; // @[Datapath.scala 81:17:@329.4]
  assign io_debug_mdr = mdr; // @[Datapath.scala 82:18:@330.4]
  assign io_debug_aluout = aluout; // @[Datapath.scala 83:21:@331.4]
  assign io_debug_pc = pc; // @[Datapath.scala 84:17:@332.4]
  assign io_debug_rd_c = regFile_io_rd_c; // @[Datapath.scala 86:19:@334.4]
  assign alu_io_A = io_ctrl_ALUSrcA ? regFile_io_rd_a : pc; // @[Datapath.scala 63:14:@304.4]
  assign alu_io_B = _T_127 ? regFile_io_rd_b : _T_126; // @[Datapath.scala 64:14:@323.4]
  assign alu_io_opcode = io_ctrl_ALUOp; // @[Datapath.scala 71:19:@324.4]
  assign regFile_clock = clock; // @[:@262.4]
  assign regFile_reset = reset; // @[:@263.4]
  assign regFile_io_ra_a = ir[25:21]; // @[Datapath.scala 54:21:@293.4]
  assign regFile_io_ra_b = ir[20:16]; // @[Datapath.scala 55:21:@295.4]
  assign regFile_io_wa = io_ctrl_RegDst ? _T_99 : _T_98; // @[Datapath.scala 56:21:@299.4]
  assign regFile_io_wd = io_ctrl_MemtoReg ? mdr : aluout; // @[Datapath.scala 57:21:@301.4]
  assign regFile_io_RegWrite = io_ctrl_RegWrite; // @[Datapath.scala 60:25:@302.4]
  assign regFile_io_ra_c = io_debug_ra_c; // @[Datapath.scala 85:21:@333.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ir = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mdr = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  aluout = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  pc = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ir <= 32'h20000000;
    end else begin
      if (io_ctrl_IRWrite) begin
        ir <= io_mem_mem_rdata;
      end
    end
    mdr <= io_mem_mem_rdata;
    aluout <= alu_io_out;
    if (reset) begin
      pc <= 32'h0;
    end else begin
      if (_T_82) begin
        if (_T_95) begin
          pc <= alu_io_out;
        end else begin
          if (_T_93) begin
            pc <= aluout;
          end else begin
            if (_T_91) begin
              pc <= _T_90;
            end else begin
              pc <= 32'h0;
            end
          end
        end
      end
    end
  end
endmodule
module Control( // @[:@336.2]
  input         clock, // @[:@337.4]
  input         reset, // @[:@338.4]
  input  [31:0] io_Inst, // @[:@339.4]
  output        io_IRWrite, // @[:@339.4]
  output        io_RegDst, // @[:@339.4]
  output        io_RegWrite, // @[:@339.4]
  output        io_ALUSrcA, // @[:@339.4]
  output [2:0]  io_ALUSrcB, // @[:@339.4]
  output [3:0]  io_ALUOp, // @[:@339.4]
  output [1:0]  io_PCSource, // @[:@339.4]
  output        io_PCWriteBEQ, // @[:@339.4]
  output        io_PCWriteBNE, // @[:@339.4]
  output        io_PCWrite, // @[:@339.4]
  output        io_IorD, // @[:@339.4]
  output        io_MemWrite, // @[:@339.4]
  output        io_MemtoReg, // @[:@339.4]
  output [3:0]  io_ctrl_dbg_cur_state, // @[:@339.4]
  output        io_ctrl_dbg_isRType, // @[:@339.4]
  output        io_ctrl_dbg_isIType, // @[:@339.4]
  output        io_ctrl_dbg_isJType, // @[:@339.4]
  output        io_ctrl_dbg_isLW, // @[:@339.4]
  output        io_ctrl_dbg_isSW, // @[:@339.4]
  output        io_ctrl_dbg_isBEQ, // @[:@339.4]
  output        io_ctrl_dbg_isBNE // @[:@339.4]
);
  wire [31:0] _T_84; // @[Control.scala 121:29:@348.4]
  wire  _T_85; // @[Control.scala 121:29:@349.4]
  wire  _T_89; // @[Control.scala 122:29:@351.4]
  wire  _T_90; // @[Control.scala 121:38:@352.4]
  wire  _T_94; // @[Control.scala 123:29:@354.4]
  wire  _T_95; // @[Control.scala 122:38:@355.4]
  wire  _T_99; // @[Control.scala 124:29:@357.4]
  wire  _T_100; // @[Control.scala 123:38:@358.4]
  wire  _T_104; // @[Control.scala 125:29:@360.4]
  wire  _T_105; // @[Control.scala 124:38:@361.4]
  wire  _T_109; // @[Control.scala 126:29:@363.4]
  wire  _T_110; // @[Control.scala 125:38:@364.4]
  wire  _T_114; // @[Control.scala 127:29:@366.4]
  wire  isRType; // @[Control.scala 126:38:@367.4]
  wire [31:0] _T_118; // @[Control.scala 128:26:@369.4]
  wire  _T_119; // @[Control.scala 128:26:@370.4]
  wire  _T_123; // @[Control.scala 129:29:@372.4]
  wire  _T_124; // @[Control.scala 128:36:@373.4]
  wire  _T_128; // @[Control.scala 130:29:@375.4]
  wire  _T_129; // @[Control.scala 129:39:@376.4]
  wire  _T_133; // @[Control.scala 131:29:@378.4]
  wire  _T_134; // @[Control.scala 130:39:@379.4]
  wire  _T_138; // @[Control.scala 132:29:@381.4]
  wire  isIType; // @[Control.scala 131:39:@382.4]
  wire  isJType; // @[Control.scala 133:25:@385.4]
  wire  isLW; // @[Control.scala 134:25:@388.4]
  wire  isSW; // @[Control.scala 135:25:@391.4]
  wire  isBEQ; // @[Control.scala 136:25:@394.4]
  wire  isBNE; // @[Control.scala 137:25:@397.4]
  reg [3:0] cur_state; // @[Control.scala 158:28:@399.4]
  reg [31:0] _RAND_0;
  wire  _T_175; // @[Conditional.scala 37:30:@414.4]
  wire  _T_181; // @[Conditional.scala 37:30:@427.6]
  wire [3:0] _T_183; // @[Mux.scala 61:16:@432.8]
  wire [3:0] _T_184; // @[Mux.scala 61:16:@433.8]
  wire [3:0] _T_185; // @[Mux.scala 61:16:@434.8]
  wire [3:0] _T_186; // @[Mux.scala 61:16:@435.8]
  wire [3:0] _T_187; // @[Mux.scala 61:16:@436.8]
  wire [3:0] _T_188; // @[Mux.scala 61:16:@437.8]
  wire [3:0] _T_189; // @[Mux.scala 61:16:@438.8]
  wire  _T_190; // @[Conditional.scala 37:30:@442.8]
  wire [3:0] _T_192; // @[Mux.scala 61:16:@447.10]
  wire [3:0] _T_193; // @[Mux.scala 61:16:@448.10]
  wire  _T_194; // @[Conditional.scala 37:30:@452.10]
  wire  _T_197; // @[Conditional.scala 37:30:@459.12]
  wire  _T_200; // @[Conditional.scala 37:30:@466.14]
  wire  _T_204; // @[Conditional.scala 37:30:@474.16]
  wire [3:0] _T_210; // @[Control.scala 84:16:@480.18]
  wire [3:0] _T_215; // @[Control.scala 84:16:@483.18]
  wire [3:0] _T_220; // @[Control.scala 84:16:@486.18]
  wire [3:0] _T_225; // @[Control.scala 84:16:@489.18]
  wire [3:0] _T_230; // @[Control.scala 84:16:@492.18]
  wire [3:0] _T_235; // @[Control.scala 84:16:@495.18]
  wire [3:0] _T_240; // @[Control.scala 84:16:@498.18]
  wire  _T_241; // @[Conditional.scala 37:30:@503.18]
  wire  _T_245; // @[Conditional.scala 37:30:@511.20]
  wire [3:0] _T_256; // @[Control.scala 84:16:@519.22]
  wire [3:0] _T_261; // @[Control.scala 84:16:@522.22]
  wire [3:0] _T_266; // @[Control.scala 84:16:@525.22]
  wire [3:0] _T_271; // @[Control.scala 84:16:@528.22]
  wire [3:0] _T_276; // @[Control.scala 84:16:@532.22]
  wire [3:0] _T_281; // @[Control.scala 84:16:@535.22]
  wire [3:0] _T_286; // @[Control.scala 84:16:@538.22]
  wire [3:0] _T_291; // @[Control.scala 84:16:@541.22]
  wire [3:0] _T_296; // @[Control.scala 84:16:@544.22]
  wire  _T_297; // @[Conditional.scala 37:30:@549.22]
  wire  _T_301; // @[Conditional.scala 37:30:@557.24]
  wire  _T_303; // @[Conditional.scala 37:30:@568.26]
  wire  _T_305; // @[Conditional.scala 37:30:@575.28]
  wire  _T_306; // @[Conditional.scala 37:30:@580.30]
  wire [3:0] _GEN_0; // @[Conditional.scala 39:67:@581.30]
  wire [3:0] _GEN_1; // @[Conditional.scala 39:67:@576.28]
  wire [1:0] _GEN_3; // @[Conditional.scala 39:67:@569.26]
  wire [3:0] _GEN_4; // @[Conditional.scala 39:67:@569.26]
  wire [3:0] _GEN_7; // @[Conditional.scala 39:67:@558.24]
  wire  _GEN_8; // @[Conditional.scala 39:67:@558.24]
  wire  _GEN_9; // @[Conditional.scala 39:67:@558.24]
  wire [1:0] _GEN_10; // @[Conditional.scala 39:67:@558.24]
  wire [3:0] _GEN_11; // @[Conditional.scala 39:67:@558.24]
  wire  _GEN_12; // @[Conditional.scala 39:67:@558.24]
  wire [3:0] _GEN_15; // @[Conditional.scala 39:67:@550.22]
  wire  _GEN_16; // @[Conditional.scala 39:67:@550.22]
  wire [3:0] _GEN_18; // @[Conditional.scala 39:67:@550.22]
  wire  _GEN_19; // @[Conditional.scala 39:67:@550.22]
  wire  _GEN_20; // @[Conditional.scala 39:67:@550.22]
  wire [1:0] _GEN_21; // @[Conditional.scala 39:67:@550.22]
  wire  _GEN_22; // @[Conditional.scala 39:67:@550.22]
  wire  _GEN_23; // @[Conditional.scala 39:67:@512.20]
  wire [3:0] _GEN_24; // @[Conditional.scala 39:67:@512.20]
  wire [3:0] _GEN_25; // @[Conditional.scala 39:67:@512.20]
  wire [3:0] _GEN_26; // @[Conditional.scala 39:67:@512.20]
  wire  _GEN_28; // @[Conditional.scala 39:67:@512.20]
  wire  _GEN_29; // @[Conditional.scala 39:67:@512.20]
  wire  _GEN_30; // @[Conditional.scala 39:67:@512.20]
  wire [1:0] _GEN_31; // @[Conditional.scala 39:67:@512.20]
  wire  _GEN_32; // @[Conditional.scala 39:67:@512.20]
  wire  _GEN_34; // @[Conditional.scala 39:67:@504.18]
  wire [3:0] _GEN_36; // @[Conditional.scala 39:67:@504.18]
  wire  _GEN_37; // @[Conditional.scala 39:67:@504.18]
  wire [3:0] _GEN_38; // @[Conditional.scala 39:67:@504.18]
  wire [3:0] _GEN_39; // @[Conditional.scala 39:67:@504.18]
  wire  _GEN_40; // @[Conditional.scala 39:67:@504.18]
  wire  _GEN_41; // @[Conditional.scala 39:67:@504.18]
  wire [1:0] _GEN_42; // @[Conditional.scala 39:67:@504.18]
  wire  _GEN_43; // @[Conditional.scala 39:67:@504.18]
  wire  _GEN_44; // @[Conditional.scala 39:67:@475.16]
  wire [3:0] _GEN_45; // @[Conditional.scala 39:67:@475.16]
  wire [3:0] _GEN_46; // @[Conditional.scala 39:67:@475.16]
  wire [3:0] _GEN_47; // @[Conditional.scala 39:67:@475.16]
  wire  _GEN_48; // @[Conditional.scala 39:67:@475.16]
  wire  _GEN_49; // @[Conditional.scala 39:67:@475.16]
  wire  _GEN_51; // @[Conditional.scala 39:67:@475.16]
  wire  _GEN_52; // @[Conditional.scala 39:67:@475.16]
  wire [1:0] _GEN_53; // @[Conditional.scala 39:67:@475.16]
  wire  _GEN_54; // @[Conditional.scala 39:67:@475.16]
  wire  _GEN_55; // @[Conditional.scala 39:67:@467.14]
  wire  _GEN_56; // @[Conditional.scala 39:67:@467.14]
  wire [3:0] _GEN_58; // @[Conditional.scala 39:67:@467.14]
  wire  _GEN_59; // @[Conditional.scala 39:67:@467.14]
  wire [3:0] _GEN_60; // @[Conditional.scala 39:67:@467.14]
  wire [3:0] _GEN_61; // @[Conditional.scala 39:67:@467.14]
  wire  _GEN_62; // @[Conditional.scala 39:67:@467.14]
  wire  _GEN_63; // @[Conditional.scala 39:67:@467.14]
  wire [1:0] _GEN_64; // @[Conditional.scala 39:67:@467.14]
  wire  _GEN_65; // @[Conditional.scala 39:67:@467.14]
  wire [3:0] _GEN_67; // @[Conditional.scala 39:67:@460.12]
  wire  _GEN_68; // @[Conditional.scala 39:67:@460.12]
  wire  _GEN_69; // @[Conditional.scala 39:67:@460.12]
  wire  _GEN_70; // @[Conditional.scala 39:67:@460.12]
  wire  _GEN_71; // @[Conditional.scala 39:67:@460.12]
  wire [3:0] _GEN_72; // @[Conditional.scala 39:67:@460.12]
  wire [3:0] _GEN_73; // @[Conditional.scala 39:67:@460.12]
  wire  _GEN_74; // @[Conditional.scala 39:67:@460.12]
  wire  _GEN_75; // @[Conditional.scala 39:67:@460.12]
  wire [1:0] _GEN_76; // @[Conditional.scala 39:67:@460.12]
  wire  _GEN_77; // @[Conditional.scala 39:67:@460.12]
  wire  _GEN_79; // @[Conditional.scala 39:67:@453.10]
  wire [3:0] _GEN_80; // @[Conditional.scala 39:67:@453.10]
  wire  _GEN_81; // @[Conditional.scala 39:67:@453.10]
  wire  _GEN_82; // @[Conditional.scala 39:67:@453.10]
  wire  _GEN_83; // @[Conditional.scala 39:67:@453.10]
  wire  _GEN_84; // @[Conditional.scala 39:67:@453.10]
  wire  _GEN_85; // @[Conditional.scala 39:67:@453.10]
  wire [3:0] _GEN_86; // @[Conditional.scala 39:67:@453.10]
  wire [3:0] _GEN_87; // @[Conditional.scala 39:67:@453.10]
  wire  _GEN_88; // @[Conditional.scala 39:67:@453.10]
  wire  _GEN_89; // @[Conditional.scala 39:67:@453.10]
  wire [1:0] _GEN_90; // @[Conditional.scala 39:67:@453.10]
  wire  _GEN_91; // @[Conditional.scala 39:67:@453.10]
  wire  _GEN_92; // @[Conditional.scala 39:67:@443.8]
  wire [3:0] _GEN_93; // @[Conditional.scala 39:67:@443.8]
  wire [3:0] _GEN_94; // @[Conditional.scala 39:67:@443.8]
  wire [3:0] _GEN_95; // @[Conditional.scala 39:67:@443.8]
  wire  _GEN_97; // @[Conditional.scala 39:67:@443.8]
  wire  _GEN_98; // @[Conditional.scala 39:67:@443.8]
  wire  _GEN_99; // @[Conditional.scala 39:67:@443.8]
  wire  _GEN_100; // @[Conditional.scala 39:67:@443.8]
  wire  _GEN_101; // @[Conditional.scala 39:67:@443.8]
  wire  _GEN_102; // @[Conditional.scala 39:67:@443.8]
  wire  _GEN_103; // @[Conditional.scala 39:67:@443.8]
  wire [1:0] _GEN_104; // @[Conditional.scala 39:67:@443.8]
  wire  _GEN_105; // @[Conditional.scala 39:67:@443.8]
  wire  _GEN_106; // @[Conditional.scala 39:67:@428.6]
  wire [3:0] _GEN_107; // @[Conditional.scala 39:67:@428.6]
  wire [3:0] _GEN_108; // @[Conditional.scala 39:67:@428.6]
  wire [3:0] _GEN_109; // @[Conditional.scala 39:67:@428.6]
  wire  _GEN_111; // @[Conditional.scala 39:67:@428.6]
  wire  _GEN_112; // @[Conditional.scala 39:67:@428.6]
  wire  _GEN_113; // @[Conditional.scala 39:67:@428.6]
  wire  _GEN_114; // @[Conditional.scala 39:67:@428.6]
  wire  _GEN_115; // @[Conditional.scala 39:67:@428.6]
  wire  _GEN_116; // @[Conditional.scala 39:67:@428.6]
  wire  _GEN_117; // @[Conditional.scala 39:67:@428.6]
  wire [1:0] _GEN_118; // @[Conditional.scala 39:67:@428.6]
  wire  _GEN_119; // @[Conditional.scala 39:67:@428.6]
  wire [3:0] _GEN_124; // @[Conditional.scala 40:58:@415.4]
  wire [3:0] _GEN_128; // @[Conditional.scala 40:58:@415.4]
  assign _T_84 = io_Inst & 32'hfc0007ff; // @[Control.scala 121:29:@348.4]
  assign _T_85 = 32'h20 == _T_84; // @[Control.scala 121:29:@349.4]
  assign _T_89 = 32'h24 == _T_84; // @[Control.scala 122:29:@351.4]
  assign _T_90 = _T_85 | _T_89; // @[Control.scala 121:38:@352.4]
  assign _T_94 = 32'h22 == _T_84; // @[Control.scala 123:29:@354.4]
  assign _T_95 = _T_90 | _T_94; // @[Control.scala 122:38:@355.4]
  assign _T_99 = 32'h25 == _T_84; // @[Control.scala 124:29:@357.4]
  assign _T_100 = _T_95 | _T_99; // @[Control.scala 123:38:@358.4]
  assign _T_104 = 32'h27 == _T_84; // @[Control.scala 125:29:@360.4]
  assign _T_105 = _T_100 | _T_104; // @[Control.scala 124:38:@361.4]
  assign _T_109 = 32'h26 == _T_84; // @[Control.scala 126:29:@363.4]
  assign _T_110 = _T_105 | _T_109; // @[Control.scala 125:38:@364.4]
  assign _T_114 = 32'h2a == _T_84; // @[Control.scala 127:29:@366.4]
  assign isRType = _T_110 | _T_114; // @[Control.scala 126:38:@367.4]
  assign _T_118 = io_Inst & 32'hfc000000; // @[Control.scala 128:26:@369.4]
  assign _T_119 = 32'h20000000 == _T_118; // @[Control.scala 128:26:@370.4]
  assign _T_123 = 32'h30000000 == _T_118; // @[Control.scala 129:29:@372.4]
  assign _T_124 = _T_119 | _T_123; // @[Control.scala 128:36:@373.4]
  assign _T_128 = 32'h34000000 == _T_118; // @[Control.scala 130:29:@375.4]
  assign _T_129 = _T_124 | _T_128; // @[Control.scala 129:39:@376.4]
  assign _T_133 = 32'h38000000 == _T_118; // @[Control.scala 131:29:@378.4]
  assign _T_134 = _T_129 | _T_133; // @[Control.scala 130:39:@379.4]
  assign _T_138 = 32'h28000000 == _T_118; // @[Control.scala 132:29:@381.4]
  assign isIType = _T_134 | _T_138; // @[Control.scala 131:39:@382.4]
  assign isJType = 32'h8000000 == _T_118; // @[Control.scala 133:25:@385.4]
  assign isLW = 32'h8c000000 == _T_118; // @[Control.scala 134:25:@388.4]
  assign isSW = 32'hac000000 == _T_118; // @[Control.scala 135:25:@391.4]
  assign isBEQ = 32'h10000000 == _T_118; // @[Control.scala 136:25:@394.4]
  assign isBNE = 32'h14000000 == _T_118; // @[Control.scala 137:25:@397.4]
  assign _T_175 = 4'h0 == cur_state; // @[Conditional.scala 37:30:@414.4]
  assign _T_181 = 4'h1 == cur_state; // @[Conditional.scala 37:30:@427.6]
  assign _T_183 = isBNE ? 4'ha : 4'hc; // @[Mux.scala 61:16:@432.8]
  assign _T_184 = isBEQ ? 4'ha : _T_183; // @[Mux.scala 61:16:@433.8]
  assign _T_185 = isSW ? 4'h2 : _T_184; // @[Mux.scala 61:16:@434.8]
  assign _T_186 = isLW ? 4'h2 : _T_185; // @[Mux.scala 61:16:@435.8]
  assign _T_187 = isJType ? 4'hb : _T_186; // @[Mux.scala 61:16:@436.8]
  assign _T_188 = isIType ? 4'h8 : _T_187; // @[Mux.scala 61:16:@437.8]
  assign _T_189 = isRType ? 4'h6 : _T_188; // @[Mux.scala 61:16:@438.8]
  assign _T_190 = 4'h2 == cur_state; // @[Conditional.scala 37:30:@442.8]
  assign _T_192 = isSW ? 4'h4 : 4'hc; // @[Mux.scala 61:16:@447.10]
  assign _T_193 = isLW ? 4'h3 : _T_192; // @[Mux.scala 61:16:@448.10]
  assign _T_194 = 4'h3 == cur_state; // @[Conditional.scala 37:30:@452.10]
  assign _T_197 = 4'h4 == cur_state; // @[Conditional.scala 37:30:@459.12]
  assign _T_200 = 4'h5 == cur_state; // @[Conditional.scala 37:30:@466.14]
  assign _T_204 = 4'h6 == cur_state; // @[Conditional.scala 37:30:@474.16]
  assign _T_210 = _T_114 ? 4'h5 : 4'hf; // @[Control.scala 84:16:@480.18]
  assign _T_215 = _T_109 ? 4'h4 : _T_210; // @[Control.scala 84:16:@483.18]
  assign _T_220 = _T_104 ? 4'hc : _T_215; // @[Control.scala 84:16:@486.18]
  assign _T_225 = _T_99 ? 4'h3 : _T_220; // @[Control.scala 84:16:@489.18]
  assign _T_230 = _T_94 ? 4'h1 : _T_225; // @[Control.scala 84:16:@492.18]
  assign _T_235 = _T_89 ? 4'h2 : _T_230; // @[Control.scala 84:16:@495.18]
  assign _T_240 = _T_85 ? 4'h0 : _T_235; // @[Control.scala 84:16:@498.18]
  assign _T_241 = 4'h7 == cur_state; // @[Conditional.scala 37:30:@503.18]
  assign _T_245 = 4'h8 == cur_state; // @[Conditional.scala 37:30:@511.20]
  assign _T_256 = _T_133 ? 4'h4 : 4'h2; // @[Control.scala 84:16:@519.22]
  assign _T_261 = _T_128 ? 4'h4 : _T_256; // @[Control.scala 84:16:@522.22]
  assign _T_266 = _T_123 ? 4'h4 : _T_261; // @[Control.scala 84:16:@525.22]
  assign _T_271 = _T_119 ? 4'h2 : _T_266; // @[Control.scala 84:16:@528.22]
  assign _T_276 = _T_138 ? 4'h5 : 4'hf; // @[Control.scala 84:16:@532.22]
  assign _T_281 = _T_133 ? 4'h4 : _T_276; // @[Control.scala 84:16:@535.22]
  assign _T_286 = _T_128 ? 4'h3 : _T_281; // @[Control.scala 84:16:@538.22]
  assign _T_291 = _T_123 ? 4'h2 : _T_286; // @[Control.scala 84:16:@541.22]
  assign _T_296 = _T_119 ? 4'h0 : _T_291; // @[Control.scala 84:16:@544.22]
  assign _T_297 = 4'h9 == cur_state; // @[Conditional.scala 37:30:@549.22]
  assign _T_301 = 4'ha == cur_state; // @[Conditional.scala 37:30:@557.24]
  assign _T_303 = 4'hb == cur_state; // @[Conditional.scala 37:30:@568.26]
  assign _T_305 = 4'hc == cur_state; // @[Conditional.scala 37:30:@575.28]
  assign _T_306 = 4'hd == cur_state; // @[Conditional.scala 37:30:@580.30]
  assign _GEN_0 = _T_306 ? 4'h0 : cur_state; // @[Conditional.scala 39:67:@581.30]
  assign _GEN_1 = _T_305 ? 4'hc : _GEN_0; // @[Conditional.scala 39:67:@576.28]
  assign _GEN_3 = _T_303 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67:@569.26]
  assign _GEN_4 = _T_303 ? 4'h0 : _GEN_1; // @[Conditional.scala 39:67:@569.26]
  assign _GEN_7 = _T_301 ? 4'h1 : 4'h0; // @[Conditional.scala 39:67:@558.24]
  assign _GEN_8 = _T_301 ? isBEQ : 1'h0; // @[Conditional.scala 39:67:@558.24]
  assign _GEN_9 = _T_301 ? isBNE : 1'h0; // @[Conditional.scala 39:67:@558.24]
  assign _GEN_10 = _T_301 ? 2'h1 : _GEN_3; // @[Conditional.scala 39:67:@558.24]
  assign _GEN_11 = _T_301 ? 4'h0 : _GEN_4; // @[Conditional.scala 39:67:@558.24]
  assign _GEN_12 = _T_301 ? 1'h0 : _T_303; // @[Conditional.scala 39:67:@558.24]
  assign _GEN_15 = _T_297 ? 4'h0 : _GEN_11; // @[Conditional.scala 39:67:@550.22]
  assign _GEN_16 = _T_297 ? 1'h0 : _T_301; // @[Conditional.scala 39:67:@550.22]
  assign _GEN_18 = _T_297 ? 4'h0 : _GEN_7; // @[Conditional.scala 39:67:@550.22]
  assign _GEN_19 = _T_297 ? 1'h0 : _GEN_8; // @[Conditional.scala 39:67:@550.22]
  assign _GEN_20 = _T_297 ? 1'h0 : _GEN_9; // @[Conditional.scala 39:67:@550.22]
  assign _GEN_21 = _T_297 ? 2'h0 : _GEN_10; // @[Conditional.scala 39:67:@550.22]
  assign _GEN_22 = _T_297 ? 1'h0 : _GEN_12; // @[Conditional.scala 39:67:@550.22]
  assign _GEN_23 = _T_245 ? 1'h1 : _GEN_16; // @[Conditional.scala 39:67:@512.20]
  assign _GEN_24 = _T_245 ? _T_271 : 4'h0; // @[Conditional.scala 39:67:@512.20]
  assign _GEN_25 = _T_245 ? _T_296 : _GEN_18; // @[Conditional.scala 39:67:@512.20]
  assign _GEN_26 = _T_245 ? 4'h9 : _GEN_15; // @[Conditional.scala 39:67:@512.20]
  assign _GEN_28 = _T_245 ? 1'h0 : _T_297; // @[Conditional.scala 39:67:@512.20]
  assign _GEN_29 = _T_245 ? 1'h0 : _GEN_19; // @[Conditional.scala 39:67:@512.20]
  assign _GEN_30 = _T_245 ? 1'h0 : _GEN_20; // @[Conditional.scala 39:67:@512.20]
  assign _GEN_31 = _T_245 ? 2'h0 : _GEN_21; // @[Conditional.scala 39:67:@512.20]
  assign _GEN_32 = _T_245 ? 1'h0 : _GEN_22; // @[Conditional.scala 39:67:@512.20]
  assign _GEN_34 = _T_241 ? 1'h1 : _GEN_28; // @[Conditional.scala 39:67:@504.18]
  assign _GEN_36 = _T_241 ? 4'h0 : _GEN_26; // @[Conditional.scala 39:67:@504.18]
  assign _GEN_37 = _T_241 ? 1'h0 : _GEN_23; // @[Conditional.scala 39:67:@504.18]
  assign _GEN_38 = _T_241 ? 4'h0 : _GEN_24; // @[Conditional.scala 39:67:@504.18]
  assign _GEN_39 = _T_241 ? 4'h0 : _GEN_25; // @[Conditional.scala 39:67:@504.18]
  assign _GEN_40 = _T_241 ? 1'h0 : _GEN_29; // @[Conditional.scala 39:67:@504.18]
  assign _GEN_41 = _T_241 ? 1'h0 : _GEN_30; // @[Conditional.scala 39:67:@504.18]
  assign _GEN_42 = _T_241 ? 2'h0 : _GEN_31; // @[Conditional.scala 39:67:@504.18]
  assign _GEN_43 = _T_241 ? 1'h0 : _GEN_32; // @[Conditional.scala 39:67:@504.18]
  assign _GEN_44 = _T_204 ? 1'h1 : _GEN_37; // @[Conditional.scala 39:67:@475.16]
  assign _GEN_45 = _T_204 ? 4'h0 : _GEN_38; // @[Conditional.scala 39:67:@475.16]
  assign _GEN_46 = _T_204 ? _T_240 : _GEN_39; // @[Conditional.scala 39:67:@475.16]
  assign _GEN_47 = _T_204 ? 4'h7 : _GEN_36; // @[Conditional.scala 39:67:@475.16]
  assign _GEN_48 = _T_204 ? 1'h0 : _T_241; // @[Conditional.scala 39:67:@475.16]
  assign _GEN_49 = _T_204 ? 1'h0 : _GEN_34; // @[Conditional.scala 39:67:@475.16]
  assign _GEN_51 = _T_204 ? 1'h0 : _GEN_40; // @[Conditional.scala 39:67:@475.16]
  assign _GEN_52 = _T_204 ? 1'h0 : _GEN_41; // @[Conditional.scala 39:67:@475.16]
  assign _GEN_53 = _T_204 ? 2'h0 : _GEN_42; // @[Conditional.scala 39:67:@475.16]
  assign _GEN_54 = _T_204 ? 1'h0 : _GEN_43; // @[Conditional.scala 39:67:@475.16]
  assign _GEN_55 = _T_200 ? 1'h0 : _GEN_48; // @[Conditional.scala 39:67:@467.14]
  assign _GEN_56 = _T_200 ? 1'h1 : _GEN_49; // @[Conditional.scala 39:67:@467.14]
  assign _GEN_58 = _T_200 ? 4'h0 : _GEN_47; // @[Conditional.scala 39:67:@467.14]
  assign _GEN_59 = _T_200 ? 1'h0 : _GEN_44; // @[Conditional.scala 39:67:@467.14]
  assign _GEN_60 = _T_200 ? 4'h0 : _GEN_45; // @[Conditional.scala 39:67:@467.14]
  assign _GEN_61 = _T_200 ? 4'h0 : _GEN_46; // @[Conditional.scala 39:67:@467.14]
  assign _GEN_62 = _T_200 ? 1'h0 : _GEN_51; // @[Conditional.scala 39:67:@467.14]
  assign _GEN_63 = _T_200 ? 1'h0 : _GEN_52; // @[Conditional.scala 39:67:@467.14]
  assign _GEN_64 = _T_200 ? 2'h0 : _GEN_53; // @[Conditional.scala 39:67:@467.14]
  assign _GEN_65 = _T_200 ? 1'h0 : _GEN_54; // @[Conditional.scala 39:67:@467.14]
  assign _GEN_67 = _T_197 ? 4'h0 : _GEN_58; // @[Conditional.scala 39:67:@460.12]
  assign _GEN_68 = _T_197 ? 1'h0 : _GEN_55; // @[Conditional.scala 39:67:@460.12]
  assign _GEN_69 = _T_197 ? 1'h0 : _GEN_56; // @[Conditional.scala 39:67:@460.12]
  assign _GEN_70 = _T_197 ? 1'h0 : _T_200; // @[Conditional.scala 39:67:@460.12]
  assign _GEN_71 = _T_197 ? 1'h0 : _GEN_59; // @[Conditional.scala 39:67:@460.12]
  assign _GEN_72 = _T_197 ? 4'h0 : _GEN_60; // @[Conditional.scala 39:67:@460.12]
  assign _GEN_73 = _T_197 ? 4'h0 : _GEN_61; // @[Conditional.scala 39:67:@460.12]
  assign _GEN_74 = _T_197 ? 1'h0 : _GEN_62; // @[Conditional.scala 39:67:@460.12]
  assign _GEN_75 = _T_197 ? 1'h0 : _GEN_63; // @[Conditional.scala 39:67:@460.12]
  assign _GEN_76 = _T_197 ? 2'h0 : _GEN_64; // @[Conditional.scala 39:67:@460.12]
  assign _GEN_77 = _T_197 ? 1'h0 : _GEN_65; // @[Conditional.scala 39:67:@460.12]
  assign _GEN_79 = _T_194 ? 1'h1 : _T_197; // @[Conditional.scala 39:67:@453.10]
  assign _GEN_80 = _T_194 ? 4'h5 : _GEN_67; // @[Conditional.scala 39:67:@453.10]
  assign _GEN_81 = _T_194 ? 1'h0 : _T_197; // @[Conditional.scala 39:67:@453.10]
  assign _GEN_82 = _T_194 ? 1'h0 : _GEN_68; // @[Conditional.scala 39:67:@453.10]
  assign _GEN_83 = _T_194 ? 1'h0 : _GEN_69; // @[Conditional.scala 39:67:@453.10]
  assign _GEN_84 = _T_194 ? 1'h0 : _GEN_70; // @[Conditional.scala 39:67:@453.10]
  assign _GEN_85 = _T_194 ? 1'h0 : _GEN_71; // @[Conditional.scala 39:67:@453.10]
  assign _GEN_86 = _T_194 ? 4'h0 : _GEN_72; // @[Conditional.scala 39:67:@453.10]
  assign _GEN_87 = _T_194 ? 4'h0 : _GEN_73; // @[Conditional.scala 39:67:@453.10]
  assign _GEN_88 = _T_194 ? 1'h0 : _GEN_74; // @[Conditional.scala 39:67:@453.10]
  assign _GEN_89 = _T_194 ? 1'h0 : _GEN_75; // @[Conditional.scala 39:67:@453.10]
  assign _GEN_90 = _T_194 ? 2'h0 : _GEN_76; // @[Conditional.scala 39:67:@453.10]
  assign _GEN_91 = _T_194 ? 1'h0 : _GEN_77; // @[Conditional.scala 39:67:@453.10]
  assign _GEN_92 = _T_190 ? 1'h1 : _GEN_85; // @[Conditional.scala 39:67:@443.8]
  assign _GEN_93 = _T_190 ? 4'h2 : _GEN_86; // @[Conditional.scala 39:67:@443.8]
  assign _GEN_94 = _T_190 ? 4'h0 : _GEN_87; // @[Conditional.scala 39:67:@443.8]
  assign _GEN_95 = _T_190 ? _T_193 : _GEN_80; // @[Conditional.scala 39:67:@443.8]
  assign _GEN_97 = _T_190 ? 1'h0 : _GEN_79; // @[Conditional.scala 39:67:@443.8]
  assign _GEN_98 = _T_190 ? 1'h0 : _GEN_81; // @[Conditional.scala 39:67:@443.8]
  assign _GEN_99 = _T_190 ? 1'h0 : _GEN_82; // @[Conditional.scala 39:67:@443.8]
  assign _GEN_100 = _T_190 ? 1'h0 : _GEN_83; // @[Conditional.scala 39:67:@443.8]
  assign _GEN_101 = _T_190 ? 1'h0 : _GEN_84; // @[Conditional.scala 39:67:@443.8]
  assign _GEN_102 = _T_190 ? 1'h0 : _GEN_88; // @[Conditional.scala 39:67:@443.8]
  assign _GEN_103 = _T_190 ? 1'h0 : _GEN_89; // @[Conditional.scala 39:67:@443.8]
  assign _GEN_104 = _T_190 ? 2'h0 : _GEN_90; // @[Conditional.scala 39:67:@443.8]
  assign _GEN_105 = _T_190 ? 1'h0 : _GEN_91; // @[Conditional.scala 39:67:@443.8]
  assign _GEN_106 = _T_181 ? 1'h1 : _GEN_92; // @[Conditional.scala 39:67:@428.6]
  assign _GEN_107 = _T_181 ? 4'h3 : _GEN_93; // @[Conditional.scala 39:67:@428.6]
  assign _GEN_108 = _T_181 ? 4'h0 : _GEN_94; // @[Conditional.scala 39:67:@428.6]
  assign _GEN_109 = _T_181 ? _T_189 : _GEN_95; // @[Conditional.scala 39:67:@428.6]
  assign _GEN_111 = _T_181 ? 1'h0 : _GEN_97; // @[Conditional.scala 39:67:@428.6]
  assign _GEN_112 = _T_181 ? 1'h0 : _GEN_98; // @[Conditional.scala 39:67:@428.6]
  assign _GEN_113 = _T_181 ? 1'h0 : _GEN_99; // @[Conditional.scala 39:67:@428.6]
  assign _GEN_114 = _T_181 ? 1'h0 : _GEN_100; // @[Conditional.scala 39:67:@428.6]
  assign _GEN_115 = _T_181 ? 1'h0 : _GEN_101; // @[Conditional.scala 39:67:@428.6]
  assign _GEN_116 = _T_181 ? 1'h0 : _GEN_102; // @[Conditional.scala 39:67:@428.6]
  assign _GEN_117 = _T_181 ? 1'h0 : _GEN_103; // @[Conditional.scala 39:67:@428.6]
  assign _GEN_118 = _T_181 ? 2'h0 : _GEN_104; // @[Conditional.scala 39:67:@428.6]
  assign _GEN_119 = _T_181 ? 1'h0 : _GEN_105; // @[Conditional.scala 39:67:@428.6]
  assign _GEN_124 = _T_175 ? 4'h1 : _GEN_107; // @[Conditional.scala 40:58:@415.4]
  assign _GEN_128 = _T_175 ? 4'h1 : _GEN_109; // @[Conditional.scala 40:58:@415.4]
  assign io_IRWrite = 4'h0 == cur_state; // @[Control.scala 140:25:@400.4 Control.scala 168:26:@419.6]
  assign io_RegDst = _T_175 ? 1'h0 : _GEN_113; // @[Control.scala 141:25:@401.4 Control.scala 219:26:@468.16 Control.scala 243:26:@505.20 Control.scala 271:25:@551.24]
  assign io_RegWrite = _T_175 ? 1'h0 : _GEN_114; // @[Control.scala 142:25:@402.4 Control.scala 220:26:@469.16 Control.scala 244:26:@506.20 Control.scala 272:26:@552.24]
  assign io_ALUSrcA = _T_175 ? 1'h0 : _GEN_106; // @[Control.scala 143:25:@403.4 Control.scala 166:26:@417.6 Control.scala 178:26:@429.8 Control.scala 194:26:@444.10 Control.scala 227:26:@476.18 Control.scala 251:26:@513.22 Control.scala 279:27:@559.26]
  assign io_ALUSrcB = _GEN_124[2:0]; // @[Control.scala 144:25:@404.4 Control.scala 169:26:@420.6 Control.scala 179:26:@430.8 Control.scala 195:26:@445.10 Control.scala 228:26:@477.18 Control.scala 252:26:@529.22 Control.scala 280:27:@560.26]
  assign io_ALUOp = _T_175 ? 4'h0 : _GEN_108; // @[Control.scala 145:25:@405.4 Control.scala 170:26:@421.6 Control.scala 180:26:@431.8 Control.scala 196:26:@446.10 Control.scala 229:26:@499.18 Control.scala 259:26:@545.22 Control.scala 281:27:@561.26]
  assign io_PCSource = _T_175 ? 2'h0 : _GEN_118; // @[Control.scala 146:25:@406.4 Control.scala 172:26:@423.6 Control.scala 284:27:@564.26 Control.scala 291:26:@571.28]
  assign io_PCWriteBEQ = _T_175 ? 1'h0 : _GEN_116; // @[Control.scala 147:25:@407.4 Control.scala 282:27:@562.26]
  assign io_PCWriteBNE = _T_175 ? 1'h0 : _GEN_117; // @[Control.scala 148:25:@408.4 Control.scala 283:27:@563.26]
  assign io_PCWrite = _T_175 ? 1'h1 : _GEN_119; // @[Control.scala 149:25:@409.4 Control.scala 171:26:@422.6 Control.scala 290:26:@570.28]
  assign io_IorD = _T_175 ? 1'h0 : _GEN_111; // @[Control.scala 150:25:@410.4 Control.scala 167:26:@418.6 Control.scala 206:26:@455.12 Control.scala 213:26:@462.14]
  assign io_MemWrite = _T_175 ? 1'h0 : _GEN_112; // @[Control.scala 152:25:@412.4 Control.scala 212:26:@461.14]
  assign io_MemtoReg = _T_175 ? 1'h0 : _GEN_115; // @[Control.scala 153:25:@413.4 Control.scala 221:26:@470.16 Control.scala 245:26:@507.20 Control.scala 273:26:@553.24]
  assign io_ctrl_dbg_cur_state = cur_state; // @[Control.scala 307:27:@584.4]
  assign io_ctrl_dbg_isRType = _T_110 | _T_114; // @[Control.scala 308:27:@585.4]
  assign io_ctrl_dbg_isIType = _T_134 | _T_138; // @[Control.scala 309:27:@586.4]
  assign io_ctrl_dbg_isJType = 32'h8000000 == _T_118; // @[Control.scala 310:27:@587.4]
  assign io_ctrl_dbg_isLW = 32'h8c000000 == _T_118; // @[Control.scala 311:27:@588.4]
  assign io_ctrl_dbg_isSW = 32'hac000000 == _T_118; // @[Control.scala 312:27:@589.4]
  assign io_ctrl_dbg_isBEQ = 32'h10000000 == _T_118; // @[Control.scala 313:27:@590.4]
  assign io_ctrl_dbg_isBNE = 32'h14000000 == _T_118; // @[Control.scala 314:27:@591.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cur_state = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cur_state <= 4'hd;
    end else begin
      if (_T_175) begin
        cur_state <= 4'h1;
      end else begin
        if (_T_181) begin
          if (isRType) begin
            cur_state <= 4'h6;
          end else begin
            if (isIType) begin
              cur_state <= 4'h8;
            end else begin
              if (isJType) begin
                cur_state <= 4'hb;
              end else begin
                if (isLW) begin
                  cur_state <= 4'h2;
                end else begin
                  if (isSW) begin
                    cur_state <= 4'h2;
                  end else begin
                    if (isBEQ) begin
                      cur_state <= 4'ha;
                    end else begin
                      if (isBNE) begin
                        cur_state <= 4'ha;
                      end else begin
                        cur_state <= 4'hc;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_190) begin
            if (isLW) begin
              cur_state <= 4'h3;
            end else begin
              if (isSW) begin
                cur_state <= 4'h4;
              end else begin
                cur_state <= 4'hc;
              end
            end
          end else begin
            if (_T_194) begin
              cur_state <= 4'h5;
            end else begin
              if (_T_197) begin
                cur_state <= 4'h0;
              end else begin
                if (_T_200) begin
                  cur_state <= 4'h0;
                end else begin
                  if (_T_204) begin
                    cur_state <= 4'h7;
                  end else begin
                    if (_T_241) begin
                      cur_state <= 4'h0;
                    end else begin
                      if (_T_245) begin
                        cur_state <= 4'h9;
                      end else begin
                        if (_T_297) begin
                          cur_state <= 4'h0;
                        end else begin
                          if (_T_301) begin
                            cur_state <= 4'h0;
                          end else begin
                            if (_T_303) begin
                              cur_state <= 4'h0;
                            end else begin
                              if (_T_305) begin
                                cur_state <= 4'hc;
                              end else begin
                                if (_T_306) begin
                                  cur_state <= 4'h0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module Mem( // @[:@593.2]
  input         clock, // @[:@594.4]
  input         reset, // @[:@595.4]
  output [31:0] io_mem_rdata, // @[:@596.4]
  input  [31:0] io_mem_addr, // @[:@596.4]
  input  [31:0] io_mem_wdata, // @[:@596.4]
  input         io_mem_wen // @[:@596.4]
);
  reg [31:0] memory_0; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_0;
  reg [31:0] memory_1; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_1;
  reg [31:0] memory_2; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_2;
  reg [31:0] memory_3; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_3;
  reg [31:0] memory_4; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_4;
  reg [31:0] memory_5; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_5;
  reg [31:0] memory_6; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_6;
  reg [31:0] memory_7; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_7;
  reg [31:0] memory_8; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_8;
  reg [31:0] memory_9; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_9;
  reg [31:0] memory_10; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_10;
  reg [31:0] memory_11; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_11;
  reg [31:0] memory_12; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_12;
  reg [31:0] memory_13; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_13;
  reg [31:0] memory_14; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_14;
  reg [31:0] memory_15; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_15;
  reg [31:0] memory_16; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_16;
  reg [31:0] memory_17; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_17;
  reg [31:0] memory_18; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_18;
  reg [31:0] memory_19; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_19;
  reg [31:0] memory_20; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_20;
  reg [31:0] memory_21; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_21;
  reg [31:0] memory_22; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_22;
  reg [31:0] memory_23; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_23;
  reg [31:0] memory_24; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_24;
  reg [31:0] memory_25; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_25;
  reg [31:0] memory_26; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_26;
  reg [31:0] memory_27; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_27;
  reg [31:0] memory_28; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_28;
  reg [31:0] memory_29; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_29;
  reg [31:0] memory_30; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_30;
  reg [31:0] memory_31; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_31;
  reg [31:0] memory_32; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_32;
  reg [31:0] memory_33; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_33;
  reg [31:0] memory_34; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_34;
  reg [31:0] memory_35; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_35;
  reg [31:0] memory_36; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_36;
  reg [31:0] memory_37; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_37;
  reg [31:0] memory_38; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_38;
  reg [31:0] memory_39; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_39;
  reg [31:0] memory_40; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_40;
  reg [31:0] memory_41; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_41;
  reg [31:0] memory_42; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_42;
  reg [31:0] memory_43; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_43;
  reg [31:0] memory_44; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_44;
  reg [31:0] memory_45; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_45;
  reg [31:0] memory_46; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_46;
  reg [31:0] memory_47; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_47;
  reg [31:0] memory_48; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_48;
  reg [31:0] memory_49; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_49;
  reg [31:0] memory_50; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_50;
  reg [31:0] memory_51; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_51;
  reg [31:0] memory_52; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_52;
  reg [31:0] memory_53; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_53;
  reg [31:0] memory_54; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_54;
  reg [31:0] memory_55; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_55;
  reg [31:0] memory_56; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_56;
  reg [31:0] memory_57; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_57;
  reg [31:0] memory_58; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_58;
  reg [31:0] memory_59; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_59;
  reg [31:0] memory_60; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_60;
  reg [31:0] memory_61; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_61;
  reg [31:0] memory_62; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_62;
  reg [31:0] memory_63; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_63;
  reg [31:0] memory_64; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_64;
  reg [31:0] memory_65; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_65;
  reg [31:0] memory_66; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_66;
  reg [31:0] memory_67; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_67;
  reg [31:0] memory_68; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_68;
  reg [31:0] memory_69; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_69;
  reg [31:0] memory_70; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_70;
  reg [31:0] memory_71; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_71;
  reg [31:0] memory_72; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_72;
  reg [31:0] memory_73; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_73;
  reg [31:0] memory_74; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_74;
  reg [31:0] memory_75; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_75;
  reg [31:0] memory_76; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_76;
  reg [31:0] memory_77; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_77;
  reg [31:0] memory_78; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_78;
  reg [31:0] memory_79; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_79;
  reg [31:0] memory_80; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_80;
  reg [31:0] memory_81; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_81;
  reg [31:0] memory_82; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_82;
  reg [31:0] memory_83; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_83;
  reg [31:0] memory_84; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_84;
  reg [31:0] memory_85; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_85;
  reg [31:0] memory_86; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_86;
  reg [31:0] memory_87; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_87;
  reg [31:0] memory_88; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_88;
  reg [31:0] memory_89; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_89;
  reg [31:0] memory_90; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_90;
  reg [31:0] memory_91; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_91;
  reg [31:0] memory_92; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_92;
  reg [31:0] memory_93; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_93;
  reg [31:0] memory_94; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_94;
  reg [31:0] memory_95; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_95;
  reg [31:0] memory_96; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_96;
  reg [31:0] memory_97; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_97;
  reg [31:0] memory_98; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_98;
  reg [31:0] memory_99; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_99;
  reg [31:0] memory_100; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_100;
  reg [31:0] memory_101; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_101;
  reg [31:0] memory_102; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_102;
  reg [31:0] memory_103; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_103;
  reg [31:0] memory_104; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_104;
  reg [31:0] memory_105; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_105;
  reg [31:0] memory_106; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_106;
  reg [31:0] memory_107; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_107;
  reg [31:0] memory_108; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_108;
  reg [31:0] memory_109; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_109;
  reg [31:0] memory_110; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_110;
  reg [31:0] memory_111; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_111;
  reg [31:0] memory_112; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_112;
  reg [31:0] memory_113; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_113;
  reg [31:0] memory_114; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_114;
  reg [31:0] memory_115; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_115;
  reg [31:0] memory_116; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_116;
  reg [31:0] memory_117; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_117;
  reg [31:0] memory_118; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_118;
  reg [31:0] memory_119; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_119;
  reg [31:0] memory_120; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_120;
  reg [31:0] memory_121; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_121;
  reg [31:0] memory_122; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_122;
  reg [31:0] memory_123; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_123;
  reg [31:0] memory_124; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_124;
  reg [31:0] memory_125; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_125;
  reg [31:0] memory_126; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_126;
  reg [31:0] memory_127; // @[Mem.scala 37:25:@727.4]
  reg [31:0] _RAND_127;
  wire  _T_921; // @[Mem.scala 39:41:@728.4]
  wire  _T_922; // @[Mem.scala 39:26:@729.4]
  wire [31:0] _GEN_0; // @[Mem.scala 39:50:@730.4]
  wire [6:0] _T_926; // @[:@733.4]
  wire [31:0] _GEN_2; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_3; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_4; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_5; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_6; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_7; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_8; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_9; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_10; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_11; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_12; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_13; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_14; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_15; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_16; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_17; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_18; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_19; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_20; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_21; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_22; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_23; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_24; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_25; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_26; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_27; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_28; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_29; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_30; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_31; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_32; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_33; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_34; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_35; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_36; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_37; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_38; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_39; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_40; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_41; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_42; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_43; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_44; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_45; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_46; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_47; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_48; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_49; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_50; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_51; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_52; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_53; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_54; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_55; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_56; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_57; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_58; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_59; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_60; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_61; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_62; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_63; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_64; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_65; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_66; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_67; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_68; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_69; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_70; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_71; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_72; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_73; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_74; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_75; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_76; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_77; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_78; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_79; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_80; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_81; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_82; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_83; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_84; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_85; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_86; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_87; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_88; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_89; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_90; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_91; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_92; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_93; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_94; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_95; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_96; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_97; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_98; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_99; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_100; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_101; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_102; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_103; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_104; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_105; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_106; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_107; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_108; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_109; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_110; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_111; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_112; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_113; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_114; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_115; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_116; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_117; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_118; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_119; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_120; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_121; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_122; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_123; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_124; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_125; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_126; // @[Mem.scala 43:32:@735.4]
  wire [31:0] _GEN_127; // @[Mem.scala 43:32:@735.4]
  wire  _T_930; // @[Mem.scala 39:41:@737.4]
  wire  _T_931; // @[Mem.scala 39:26:@738.4]
  wire [31:0] _GEN_129; // @[Mem.scala 39:50:@739.4]
  wire  _T_939; // @[Mem.scala 39:41:@746.4]
  wire  _T_940; // @[Mem.scala 39:26:@747.4]
  wire [31:0] _GEN_258; // @[Mem.scala 39:50:@748.4]
  wire  _T_948; // @[Mem.scala 39:41:@755.4]
  wire  _T_949; // @[Mem.scala 39:26:@756.4]
  wire [31:0] _GEN_387; // @[Mem.scala 39:50:@757.4]
  wire  _T_957; // @[Mem.scala 39:41:@764.4]
  wire  _T_958; // @[Mem.scala 39:26:@765.4]
  wire [31:0] _GEN_516; // @[Mem.scala 39:50:@766.4]
  wire  _T_966; // @[Mem.scala 39:41:@773.4]
  wire  _T_967; // @[Mem.scala 39:26:@774.4]
  wire [31:0] _GEN_645; // @[Mem.scala 39:50:@775.4]
  wire  _T_975; // @[Mem.scala 39:41:@782.4]
  wire  _T_976; // @[Mem.scala 39:26:@783.4]
  wire [31:0] _GEN_774; // @[Mem.scala 39:50:@784.4]
  wire  _T_984; // @[Mem.scala 39:41:@791.4]
  wire  _T_985; // @[Mem.scala 39:26:@792.4]
  wire [31:0] _GEN_903; // @[Mem.scala 39:50:@793.4]
  wire  _T_993; // @[Mem.scala 39:41:@800.4]
  wire  _T_994; // @[Mem.scala 39:26:@801.4]
  wire [31:0] _GEN_1032; // @[Mem.scala 39:50:@802.4]
  wire  _T_1002; // @[Mem.scala 39:41:@809.4]
  wire  _T_1003; // @[Mem.scala 39:26:@810.4]
  wire [31:0] _GEN_1161; // @[Mem.scala 39:50:@811.4]
  wire  _T_1011; // @[Mem.scala 39:41:@818.4]
  wire  _T_1012; // @[Mem.scala 39:26:@819.4]
  wire [31:0] _GEN_1290; // @[Mem.scala 39:50:@820.4]
  wire  _T_1020; // @[Mem.scala 39:41:@827.4]
  wire  _T_1021; // @[Mem.scala 39:26:@828.4]
  wire [31:0] _GEN_1419; // @[Mem.scala 39:50:@829.4]
  wire  _T_1029; // @[Mem.scala 39:41:@836.4]
  wire  _T_1030; // @[Mem.scala 39:26:@837.4]
  wire [31:0] _GEN_1548; // @[Mem.scala 39:50:@838.4]
  wire  _T_1038; // @[Mem.scala 39:41:@845.4]
  wire  _T_1039; // @[Mem.scala 39:26:@846.4]
  wire [31:0] _GEN_1677; // @[Mem.scala 39:50:@847.4]
  wire  _T_1047; // @[Mem.scala 39:41:@854.4]
  wire  _T_1048; // @[Mem.scala 39:26:@855.4]
  wire [31:0] _GEN_1806; // @[Mem.scala 39:50:@856.4]
  wire  _T_1056; // @[Mem.scala 39:41:@863.4]
  wire  _T_1057; // @[Mem.scala 39:26:@864.4]
  wire [31:0] _GEN_1935; // @[Mem.scala 39:50:@865.4]
  wire  _T_1065; // @[Mem.scala 39:41:@872.4]
  wire  _T_1066; // @[Mem.scala 39:26:@873.4]
  wire [31:0] _GEN_2064; // @[Mem.scala 39:50:@874.4]
  wire  _T_1074; // @[Mem.scala 39:41:@881.4]
  wire  _T_1075; // @[Mem.scala 39:26:@882.4]
  wire [31:0] _GEN_2193; // @[Mem.scala 39:50:@883.4]
  wire  _T_1083; // @[Mem.scala 39:41:@890.4]
  wire  _T_1084; // @[Mem.scala 39:26:@891.4]
  wire [31:0] _GEN_2322; // @[Mem.scala 39:50:@892.4]
  wire  _T_1092; // @[Mem.scala 39:41:@899.4]
  wire  _T_1093; // @[Mem.scala 39:26:@900.4]
  wire [31:0] _GEN_2451; // @[Mem.scala 39:50:@901.4]
  wire  _T_1101; // @[Mem.scala 39:41:@908.4]
  wire  _T_1102; // @[Mem.scala 39:26:@909.4]
  wire [31:0] _GEN_2580; // @[Mem.scala 39:50:@910.4]
  wire  _T_1110; // @[Mem.scala 39:41:@917.4]
  wire  _T_1111; // @[Mem.scala 39:26:@918.4]
  wire [31:0] _GEN_2709; // @[Mem.scala 39:50:@919.4]
  wire  _T_1119; // @[Mem.scala 39:41:@926.4]
  wire  _T_1120; // @[Mem.scala 39:26:@927.4]
  wire [31:0] _GEN_2838; // @[Mem.scala 39:50:@928.4]
  wire  _T_1128; // @[Mem.scala 39:41:@935.4]
  wire  _T_1129; // @[Mem.scala 39:26:@936.4]
  wire [31:0] _GEN_2967; // @[Mem.scala 39:50:@937.4]
  wire  _T_1137; // @[Mem.scala 39:41:@944.4]
  wire  _T_1138; // @[Mem.scala 39:26:@945.4]
  wire [31:0] _GEN_3096; // @[Mem.scala 39:50:@946.4]
  wire  _T_1146; // @[Mem.scala 39:41:@953.4]
  wire  _T_1147; // @[Mem.scala 39:26:@954.4]
  wire [31:0] _GEN_3225; // @[Mem.scala 39:50:@955.4]
  wire  _T_1155; // @[Mem.scala 39:41:@962.4]
  wire  _T_1156; // @[Mem.scala 39:26:@963.4]
  wire [31:0] _GEN_3354; // @[Mem.scala 39:50:@964.4]
  wire  _T_1164; // @[Mem.scala 39:41:@971.4]
  wire  _T_1165; // @[Mem.scala 39:26:@972.4]
  wire [31:0] _GEN_3483; // @[Mem.scala 39:50:@973.4]
  wire  _T_1173; // @[Mem.scala 39:41:@980.4]
  wire  _T_1174; // @[Mem.scala 39:26:@981.4]
  wire [31:0] _GEN_3612; // @[Mem.scala 39:50:@982.4]
  wire  _T_1182; // @[Mem.scala 39:41:@989.4]
  wire  _T_1183; // @[Mem.scala 39:26:@990.4]
  wire [31:0] _GEN_3741; // @[Mem.scala 39:50:@991.4]
  wire  _T_1191; // @[Mem.scala 39:41:@998.4]
  wire  _T_1192; // @[Mem.scala 39:26:@999.4]
  wire [31:0] _GEN_3870; // @[Mem.scala 39:50:@1000.4]
  wire  _T_1200; // @[Mem.scala 39:41:@1007.4]
  wire  _T_1201; // @[Mem.scala 39:26:@1008.4]
  wire [31:0] _GEN_3999; // @[Mem.scala 39:50:@1009.4]
  wire  _T_1209; // @[Mem.scala 39:41:@1016.4]
  wire  _T_1210; // @[Mem.scala 39:26:@1017.4]
  wire [31:0] _GEN_4128; // @[Mem.scala 39:50:@1018.4]
  wire  _T_1218; // @[Mem.scala 39:41:@1025.4]
  wire  _T_1219; // @[Mem.scala 39:26:@1026.4]
  wire [31:0] _GEN_4257; // @[Mem.scala 39:50:@1027.4]
  wire  _T_1227; // @[Mem.scala 39:41:@1034.4]
  wire  _T_1228; // @[Mem.scala 39:26:@1035.4]
  wire [31:0] _GEN_4386; // @[Mem.scala 39:50:@1036.4]
  wire  _T_1236; // @[Mem.scala 39:41:@1043.4]
  wire  _T_1237; // @[Mem.scala 39:26:@1044.4]
  wire [31:0] _GEN_4515; // @[Mem.scala 39:50:@1045.4]
  wire  _T_1245; // @[Mem.scala 39:41:@1052.4]
  wire  _T_1246; // @[Mem.scala 39:26:@1053.4]
  wire [31:0] _GEN_4644; // @[Mem.scala 39:50:@1054.4]
  wire  _T_1254; // @[Mem.scala 39:41:@1061.4]
  wire  _T_1255; // @[Mem.scala 39:26:@1062.4]
  wire [31:0] _GEN_4773; // @[Mem.scala 39:50:@1063.4]
  wire  _T_1263; // @[Mem.scala 39:41:@1070.4]
  wire  _T_1264; // @[Mem.scala 39:26:@1071.4]
  wire [31:0] _GEN_4902; // @[Mem.scala 39:50:@1072.4]
  wire  _T_1272; // @[Mem.scala 39:41:@1079.4]
  wire  _T_1273; // @[Mem.scala 39:26:@1080.4]
  wire [31:0] _GEN_5031; // @[Mem.scala 39:50:@1081.4]
  wire  _T_1281; // @[Mem.scala 39:41:@1088.4]
  wire  _T_1282; // @[Mem.scala 39:26:@1089.4]
  wire [31:0] _GEN_5160; // @[Mem.scala 39:50:@1090.4]
  wire  _T_1290; // @[Mem.scala 39:41:@1097.4]
  wire  _T_1291; // @[Mem.scala 39:26:@1098.4]
  wire [31:0] _GEN_5289; // @[Mem.scala 39:50:@1099.4]
  wire  _T_1299; // @[Mem.scala 39:41:@1106.4]
  wire  _T_1300; // @[Mem.scala 39:26:@1107.4]
  wire [31:0] _GEN_5418; // @[Mem.scala 39:50:@1108.4]
  wire  _T_1308; // @[Mem.scala 39:41:@1115.4]
  wire  _T_1309; // @[Mem.scala 39:26:@1116.4]
  wire [31:0] _GEN_5547; // @[Mem.scala 39:50:@1117.4]
  wire  _T_1317; // @[Mem.scala 39:41:@1124.4]
  wire  _T_1318; // @[Mem.scala 39:26:@1125.4]
  wire [31:0] _GEN_5676; // @[Mem.scala 39:50:@1126.4]
  wire  _T_1326; // @[Mem.scala 39:41:@1133.4]
  wire  _T_1327; // @[Mem.scala 39:26:@1134.4]
  wire [31:0] _GEN_5805; // @[Mem.scala 39:50:@1135.4]
  wire  _T_1335; // @[Mem.scala 39:41:@1142.4]
  wire  _T_1336; // @[Mem.scala 39:26:@1143.4]
  wire [31:0] _GEN_5934; // @[Mem.scala 39:50:@1144.4]
  wire  _T_1344; // @[Mem.scala 39:41:@1151.4]
  wire  _T_1345; // @[Mem.scala 39:26:@1152.4]
  wire [31:0] _GEN_6063; // @[Mem.scala 39:50:@1153.4]
  wire  _T_1353; // @[Mem.scala 39:41:@1160.4]
  wire  _T_1354; // @[Mem.scala 39:26:@1161.4]
  wire [31:0] _GEN_6192; // @[Mem.scala 39:50:@1162.4]
  wire  _T_1362; // @[Mem.scala 39:41:@1169.4]
  wire  _T_1363; // @[Mem.scala 39:26:@1170.4]
  wire [31:0] _GEN_6321; // @[Mem.scala 39:50:@1171.4]
  wire  _T_1371; // @[Mem.scala 39:41:@1178.4]
  wire  _T_1372; // @[Mem.scala 39:26:@1179.4]
  wire [31:0] _GEN_6450; // @[Mem.scala 39:50:@1180.4]
  wire  _T_1380; // @[Mem.scala 39:41:@1187.4]
  wire  _T_1381; // @[Mem.scala 39:26:@1188.4]
  wire [31:0] _GEN_6579; // @[Mem.scala 39:50:@1189.4]
  wire  _T_1389; // @[Mem.scala 39:41:@1196.4]
  wire  _T_1390; // @[Mem.scala 39:26:@1197.4]
  wire [31:0] _GEN_6708; // @[Mem.scala 39:50:@1198.4]
  wire  _T_1398; // @[Mem.scala 39:41:@1205.4]
  wire  _T_1399; // @[Mem.scala 39:26:@1206.4]
  wire [31:0] _GEN_6837; // @[Mem.scala 39:50:@1207.4]
  wire  _T_1407; // @[Mem.scala 39:41:@1214.4]
  wire  _T_1408; // @[Mem.scala 39:26:@1215.4]
  wire [31:0] _GEN_6966; // @[Mem.scala 39:50:@1216.4]
  wire  _T_1416; // @[Mem.scala 39:41:@1223.4]
  wire  _T_1417; // @[Mem.scala 39:26:@1224.4]
  wire [31:0] _GEN_7095; // @[Mem.scala 39:50:@1225.4]
  wire  _T_1425; // @[Mem.scala 39:41:@1232.4]
  wire  _T_1426; // @[Mem.scala 39:26:@1233.4]
  wire [31:0] _GEN_7224; // @[Mem.scala 39:50:@1234.4]
  wire  _T_1434; // @[Mem.scala 39:41:@1241.4]
  wire  _T_1435; // @[Mem.scala 39:26:@1242.4]
  wire [31:0] _GEN_7353; // @[Mem.scala 39:50:@1243.4]
  wire  _T_1443; // @[Mem.scala 39:41:@1250.4]
  wire  _T_1444; // @[Mem.scala 39:26:@1251.4]
  wire [31:0] _GEN_7482; // @[Mem.scala 39:50:@1252.4]
  wire  _T_1452; // @[Mem.scala 39:41:@1259.4]
  wire  _T_1453; // @[Mem.scala 39:26:@1260.4]
  wire [31:0] _GEN_7611; // @[Mem.scala 39:50:@1261.4]
  wire  _T_1461; // @[Mem.scala 39:41:@1268.4]
  wire  _T_1462; // @[Mem.scala 39:26:@1269.4]
  wire [31:0] _GEN_7740; // @[Mem.scala 39:50:@1270.4]
  wire  _T_1470; // @[Mem.scala 39:41:@1277.4]
  wire  _T_1471; // @[Mem.scala 39:26:@1278.4]
  wire [31:0] _GEN_7869; // @[Mem.scala 39:50:@1279.4]
  wire  _T_1479; // @[Mem.scala 39:41:@1286.4]
  wire  _T_1480; // @[Mem.scala 39:26:@1287.4]
  wire [31:0] _GEN_7998; // @[Mem.scala 39:50:@1288.4]
  wire  _T_1488; // @[Mem.scala 39:41:@1295.4]
  wire  _T_1489; // @[Mem.scala 39:26:@1296.4]
  wire [31:0] _GEN_8127; // @[Mem.scala 39:50:@1297.4]
  wire  _T_1497; // @[Mem.scala 39:41:@1304.4]
  wire  _T_1498; // @[Mem.scala 39:26:@1305.4]
  wire [31:0] _GEN_8256; // @[Mem.scala 39:50:@1306.4]
  wire  _T_1506; // @[Mem.scala 39:41:@1313.4]
  wire  _T_1507; // @[Mem.scala 39:26:@1314.4]
  wire [31:0] _GEN_8385; // @[Mem.scala 39:50:@1315.4]
  wire  _T_1515; // @[Mem.scala 39:41:@1322.4]
  wire  _T_1516; // @[Mem.scala 39:26:@1323.4]
  wire [31:0] _GEN_8514; // @[Mem.scala 39:50:@1324.4]
  wire  _T_1524; // @[Mem.scala 39:41:@1331.4]
  wire  _T_1525; // @[Mem.scala 39:26:@1332.4]
  wire [31:0] _GEN_8643; // @[Mem.scala 39:50:@1333.4]
  wire  _T_1533; // @[Mem.scala 39:41:@1340.4]
  wire  _T_1534; // @[Mem.scala 39:26:@1341.4]
  wire [31:0] _GEN_8772; // @[Mem.scala 39:50:@1342.4]
  wire  _T_1542; // @[Mem.scala 39:41:@1349.4]
  wire  _T_1543; // @[Mem.scala 39:26:@1350.4]
  wire [31:0] _GEN_8901; // @[Mem.scala 39:50:@1351.4]
  wire  _T_1551; // @[Mem.scala 39:41:@1358.4]
  wire  _T_1552; // @[Mem.scala 39:26:@1359.4]
  wire [31:0] _GEN_9030; // @[Mem.scala 39:50:@1360.4]
  wire  _T_1560; // @[Mem.scala 39:41:@1367.4]
  wire  _T_1561; // @[Mem.scala 39:26:@1368.4]
  wire [31:0] _GEN_9159; // @[Mem.scala 39:50:@1369.4]
  wire  _T_1569; // @[Mem.scala 39:41:@1376.4]
  wire  _T_1570; // @[Mem.scala 39:26:@1377.4]
  wire [31:0] _GEN_9288; // @[Mem.scala 39:50:@1378.4]
  wire  _T_1578; // @[Mem.scala 39:41:@1385.4]
  wire  _T_1579; // @[Mem.scala 39:26:@1386.4]
  wire [31:0] _GEN_9417; // @[Mem.scala 39:50:@1387.4]
  wire  _T_1587; // @[Mem.scala 39:41:@1394.4]
  wire  _T_1588; // @[Mem.scala 39:26:@1395.4]
  wire [31:0] _GEN_9546; // @[Mem.scala 39:50:@1396.4]
  wire  _T_1596; // @[Mem.scala 39:41:@1403.4]
  wire  _T_1597; // @[Mem.scala 39:26:@1404.4]
  wire [31:0] _GEN_9675; // @[Mem.scala 39:50:@1405.4]
  wire  _T_1605; // @[Mem.scala 39:41:@1412.4]
  wire  _T_1606; // @[Mem.scala 39:26:@1413.4]
  wire [31:0] _GEN_9804; // @[Mem.scala 39:50:@1414.4]
  wire  _T_1614; // @[Mem.scala 39:41:@1421.4]
  wire  _T_1615; // @[Mem.scala 39:26:@1422.4]
  wire [31:0] _GEN_9933; // @[Mem.scala 39:50:@1423.4]
  wire  _T_1623; // @[Mem.scala 39:41:@1430.4]
  wire  _T_1624; // @[Mem.scala 39:26:@1431.4]
  wire [31:0] _GEN_10062; // @[Mem.scala 39:50:@1432.4]
  wire  _T_1632; // @[Mem.scala 39:41:@1439.4]
  wire  _T_1633; // @[Mem.scala 39:26:@1440.4]
  wire [31:0] _GEN_10191; // @[Mem.scala 39:50:@1441.4]
  wire  _T_1641; // @[Mem.scala 39:41:@1448.4]
  wire  _T_1642; // @[Mem.scala 39:26:@1449.4]
  wire [31:0] _GEN_10320; // @[Mem.scala 39:50:@1450.4]
  wire  _T_1650; // @[Mem.scala 39:41:@1457.4]
  wire  _T_1651; // @[Mem.scala 39:26:@1458.4]
  wire [31:0] _GEN_10449; // @[Mem.scala 39:50:@1459.4]
  wire  _T_1659; // @[Mem.scala 39:41:@1466.4]
  wire  _T_1660; // @[Mem.scala 39:26:@1467.4]
  wire [31:0] _GEN_10578; // @[Mem.scala 39:50:@1468.4]
  wire  _T_1668; // @[Mem.scala 39:41:@1475.4]
  wire  _T_1669; // @[Mem.scala 39:26:@1476.4]
  wire [31:0] _GEN_10707; // @[Mem.scala 39:50:@1477.4]
  wire  _T_1677; // @[Mem.scala 39:41:@1484.4]
  wire  _T_1678; // @[Mem.scala 39:26:@1485.4]
  wire [31:0] _GEN_10836; // @[Mem.scala 39:50:@1486.4]
  wire  _T_1686; // @[Mem.scala 39:41:@1493.4]
  wire  _T_1687; // @[Mem.scala 39:26:@1494.4]
  wire [31:0] _GEN_10965; // @[Mem.scala 39:50:@1495.4]
  wire  _T_1695; // @[Mem.scala 39:41:@1502.4]
  wire  _T_1696; // @[Mem.scala 39:26:@1503.4]
  wire [31:0] _GEN_11094; // @[Mem.scala 39:50:@1504.4]
  wire  _T_1704; // @[Mem.scala 39:41:@1511.4]
  wire  _T_1705; // @[Mem.scala 39:26:@1512.4]
  wire [31:0] _GEN_11223; // @[Mem.scala 39:50:@1513.4]
  wire  _T_1713; // @[Mem.scala 39:41:@1520.4]
  wire  _T_1714; // @[Mem.scala 39:26:@1521.4]
  wire [31:0] _GEN_11352; // @[Mem.scala 39:50:@1522.4]
  wire  _T_1722; // @[Mem.scala 39:41:@1529.4]
  wire  _T_1723; // @[Mem.scala 39:26:@1530.4]
  wire [31:0] _GEN_11481; // @[Mem.scala 39:50:@1531.4]
  wire  _T_1731; // @[Mem.scala 39:41:@1538.4]
  wire  _T_1732; // @[Mem.scala 39:26:@1539.4]
  wire [31:0] _GEN_11610; // @[Mem.scala 39:50:@1540.4]
  wire  _T_1740; // @[Mem.scala 39:41:@1547.4]
  wire  _T_1741; // @[Mem.scala 39:26:@1548.4]
  wire [31:0] _GEN_11739; // @[Mem.scala 39:50:@1549.4]
  wire  _T_1749; // @[Mem.scala 39:41:@1556.4]
  wire  _T_1750; // @[Mem.scala 39:26:@1557.4]
  wire [31:0] _GEN_11868; // @[Mem.scala 39:50:@1558.4]
  wire  _T_1758; // @[Mem.scala 39:41:@1565.4]
  wire  _T_1759; // @[Mem.scala 39:26:@1566.4]
  wire [31:0] _GEN_11997; // @[Mem.scala 39:50:@1567.4]
  wire  _T_1767; // @[Mem.scala 39:41:@1574.4]
  wire  _T_1768; // @[Mem.scala 39:26:@1575.4]
  wire [31:0] _GEN_12126; // @[Mem.scala 39:50:@1576.4]
  wire  _T_1776; // @[Mem.scala 39:41:@1583.4]
  wire  _T_1777; // @[Mem.scala 39:26:@1584.4]
  wire [31:0] _GEN_12255; // @[Mem.scala 39:50:@1585.4]
  wire  _T_1785; // @[Mem.scala 39:41:@1592.4]
  wire  _T_1786; // @[Mem.scala 39:26:@1593.4]
  wire [31:0] _GEN_12384; // @[Mem.scala 39:50:@1594.4]
  wire  _T_1794; // @[Mem.scala 39:41:@1601.4]
  wire  _T_1795; // @[Mem.scala 39:26:@1602.4]
  wire [31:0] _GEN_12513; // @[Mem.scala 39:50:@1603.4]
  wire  _T_1803; // @[Mem.scala 39:41:@1610.4]
  wire  _T_1804; // @[Mem.scala 39:26:@1611.4]
  wire [31:0] _GEN_12642; // @[Mem.scala 39:50:@1612.4]
  wire  _T_1812; // @[Mem.scala 39:41:@1619.4]
  wire  _T_1813; // @[Mem.scala 39:26:@1620.4]
  wire [31:0] _GEN_12771; // @[Mem.scala 39:50:@1621.4]
  wire  _T_1821; // @[Mem.scala 39:41:@1628.4]
  wire  _T_1822; // @[Mem.scala 39:26:@1629.4]
  wire [31:0] _GEN_12900; // @[Mem.scala 39:50:@1630.4]
  wire  _T_1830; // @[Mem.scala 39:41:@1637.4]
  wire  _T_1831; // @[Mem.scala 39:26:@1638.4]
  wire [31:0] _GEN_13029; // @[Mem.scala 39:50:@1639.4]
  wire  _T_1839; // @[Mem.scala 39:41:@1646.4]
  wire  _T_1840; // @[Mem.scala 39:26:@1647.4]
  wire [31:0] _GEN_13158; // @[Mem.scala 39:50:@1648.4]
  wire  _T_1848; // @[Mem.scala 39:41:@1655.4]
  wire  _T_1849; // @[Mem.scala 39:26:@1656.4]
  wire [31:0] _GEN_13287; // @[Mem.scala 39:50:@1657.4]
  wire  _T_1857; // @[Mem.scala 39:41:@1664.4]
  wire  _T_1858; // @[Mem.scala 39:26:@1665.4]
  wire [31:0] _GEN_13416; // @[Mem.scala 39:50:@1666.4]
  wire  _T_1866; // @[Mem.scala 39:41:@1673.4]
  wire  _T_1867; // @[Mem.scala 39:26:@1674.4]
  wire [31:0] _GEN_13545; // @[Mem.scala 39:50:@1675.4]
  wire  _T_1875; // @[Mem.scala 39:41:@1682.4]
  wire  _T_1876; // @[Mem.scala 39:26:@1683.4]
  wire [31:0] _GEN_13674; // @[Mem.scala 39:50:@1684.4]
  wire  _T_1884; // @[Mem.scala 39:41:@1691.4]
  wire  _T_1885; // @[Mem.scala 39:26:@1692.4]
  wire [31:0] _GEN_13803; // @[Mem.scala 39:50:@1693.4]
  wire  _T_1893; // @[Mem.scala 39:41:@1700.4]
  wire  _T_1894; // @[Mem.scala 39:26:@1701.4]
  wire [31:0] _GEN_13932; // @[Mem.scala 39:50:@1702.4]
  wire  _T_1902; // @[Mem.scala 39:41:@1709.4]
  wire  _T_1903; // @[Mem.scala 39:26:@1710.4]
  wire [31:0] _GEN_14061; // @[Mem.scala 39:50:@1711.4]
  wire  _T_1911; // @[Mem.scala 39:41:@1718.4]
  wire  _T_1912; // @[Mem.scala 39:26:@1719.4]
  wire [31:0] _GEN_14190; // @[Mem.scala 39:50:@1720.4]
  wire  _T_1920; // @[Mem.scala 39:41:@1727.4]
  wire  _T_1921; // @[Mem.scala 39:26:@1728.4]
  wire [31:0] _GEN_14319; // @[Mem.scala 39:50:@1729.4]
  wire  _T_1929; // @[Mem.scala 39:41:@1736.4]
  wire  _T_1930; // @[Mem.scala 39:26:@1737.4]
  wire [31:0] _GEN_14448; // @[Mem.scala 39:50:@1738.4]
  wire  _T_1938; // @[Mem.scala 39:41:@1745.4]
  wire  _T_1939; // @[Mem.scala 39:26:@1746.4]
  wire [31:0] _GEN_14577; // @[Mem.scala 39:50:@1747.4]
  wire  _T_1947; // @[Mem.scala 39:41:@1754.4]
  wire  _T_1948; // @[Mem.scala 39:26:@1755.4]
  wire [31:0] _GEN_14706; // @[Mem.scala 39:50:@1756.4]
  wire  _T_1956; // @[Mem.scala 39:41:@1763.4]
  wire  _T_1957; // @[Mem.scala 39:26:@1764.4]
  wire [31:0] _GEN_14835; // @[Mem.scala 39:50:@1765.4]
  wire  _T_1965; // @[Mem.scala 39:41:@1772.4]
  wire  _T_1966; // @[Mem.scala 39:26:@1773.4]
  wire [31:0] _GEN_14964; // @[Mem.scala 39:50:@1774.4]
  wire  _T_1974; // @[Mem.scala 39:41:@1781.4]
  wire  _T_1975; // @[Mem.scala 39:26:@1782.4]
  wire [31:0] _GEN_15093; // @[Mem.scala 39:50:@1783.4]
  wire  _T_1983; // @[Mem.scala 39:41:@1790.4]
  wire  _T_1984; // @[Mem.scala 39:26:@1791.4]
  wire [31:0] _GEN_15222; // @[Mem.scala 39:50:@1792.4]
  wire  _T_1992; // @[Mem.scala 39:41:@1799.4]
  wire  _T_1993; // @[Mem.scala 39:26:@1800.4]
  wire [31:0] _GEN_15351; // @[Mem.scala 39:50:@1801.4]
  wire  _T_2001; // @[Mem.scala 39:41:@1808.4]
  wire  _T_2002; // @[Mem.scala 39:26:@1809.4]
  wire [31:0] _GEN_15480; // @[Mem.scala 39:50:@1810.4]
  wire  _T_2010; // @[Mem.scala 39:41:@1817.4]
  wire  _T_2011; // @[Mem.scala 39:26:@1818.4]
  wire [31:0] _GEN_15609; // @[Mem.scala 39:50:@1819.4]
  wire  _T_2019; // @[Mem.scala 39:41:@1826.4]
  wire  _T_2020; // @[Mem.scala 39:26:@1827.4]
  wire [31:0] _GEN_15738; // @[Mem.scala 39:50:@1828.4]
  wire  _T_2028; // @[Mem.scala 39:41:@1835.4]
  wire  _T_2029; // @[Mem.scala 39:26:@1836.4]
  wire [31:0] _GEN_15867; // @[Mem.scala 39:50:@1837.4]
  wire  _T_2037; // @[Mem.scala 39:41:@1844.4]
  wire  _T_2038; // @[Mem.scala 39:26:@1845.4]
  wire [31:0] _GEN_15996; // @[Mem.scala 39:50:@1846.4]
  wire  _T_2046; // @[Mem.scala 39:41:@1853.4]
  wire  _T_2047; // @[Mem.scala 39:26:@1854.4]
  wire [31:0] _GEN_16125; // @[Mem.scala 39:50:@1855.4]
  wire  _T_2055; // @[Mem.scala 39:41:@1862.4]
  wire  _T_2056; // @[Mem.scala 39:26:@1863.4]
  wire [31:0] _GEN_16254; // @[Mem.scala 39:50:@1864.4]
  wire  _T_2064; // @[Mem.scala 39:41:@1871.4]
  wire  _T_2065; // @[Mem.scala 39:26:@1872.4]
  wire [31:0] _GEN_16383; // @[Mem.scala 39:50:@1873.4]
  reg [31:0] _T_2071; // @[Mem.scala 43:32:@1877.4]
  reg [31:0] _RAND_128;
  assign _T_921 = io_mem_addr == 32'h0; // @[Mem.scala 39:41:@728.4]
  assign _T_922 = io_mem_wen & _T_921; // @[Mem.scala 39:26:@729.4]
  assign _GEN_0 = _T_922 ? io_mem_wdata : memory_0; // @[Mem.scala 39:50:@730.4]
  assign _T_926 = io_mem_addr[6:0]; // @[:@733.4]
  assign _GEN_2 = 7'h1 == _T_926 ? memory_1 : memory_0; // @[Mem.scala 43:32:@735.4]
  assign _GEN_3 = 7'h2 == _T_926 ? memory_2 : _GEN_2; // @[Mem.scala 43:32:@735.4]
  assign _GEN_4 = 7'h3 == _T_926 ? memory_3 : _GEN_3; // @[Mem.scala 43:32:@735.4]
  assign _GEN_5 = 7'h4 == _T_926 ? memory_4 : _GEN_4; // @[Mem.scala 43:32:@735.4]
  assign _GEN_6 = 7'h5 == _T_926 ? memory_5 : _GEN_5; // @[Mem.scala 43:32:@735.4]
  assign _GEN_7 = 7'h6 == _T_926 ? memory_6 : _GEN_6; // @[Mem.scala 43:32:@735.4]
  assign _GEN_8 = 7'h7 == _T_926 ? memory_7 : _GEN_7; // @[Mem.scala 43:32:@735.4]
  assign _GEN_9 = 7'h8 == _T_926 ? memory_8 : _GEN_8; // @[Mem.scala 43:32:@735.4]
  assign _GEN_10 = 7'h9 == _T_926 ? memory_9 : _GEN_9; // @[Mem.scala 43:32:@735.4]
  assign _GEN_11 = 7'ha == _T_926 ? memory_10 : _GEN_10; // @[Mem.scala 43:32:@735.4]
  assign _GEN_12 = 7'hb == _T_926 ? memory_11 : _GEN_11; // @[Mem.scala 43:32:@735.4]
  assign _GEN_13 = 7'hc == _T_926 ? memory_12 : _GEN_12; // @[Mem.scala 43:32:@735.4]
  assign _GEN_14 = 7'hd == _T_926 ? memory_13 : _GEN_13; // @[Mem.scala 43:32:@735.4]
  assign _GEN_15 = 7'he == _T_926 ? memory_14 : _GEN_14; // @[Mem.scala 43:32:@735.4]
  assign _GEN_16 = 7'hf == _T_926 ? memory_15 : _GEN_15; // @[Mem.scala 43:32:@735.4]
  assign _GEN_17 = 7'h10 == _T_926 ? memory_16 : _GEN_16; // @[Mem.scala 43:32:@735.4]
  assign _GEN_18 = 7'h11 == _T_926 ? memory_17 : _GEN_17; // @[Mem.scala 43:32:@735.4]
  assign _GEN_19 = 7'h12 == _T_926 ? memory_18 : _GEN_18; // @[Mem.scala 43:32:@735.4]
  assign _GEN_20 = 7'h13 == _T_926 ? memory_19 : _GEN_19; // @[Mem.scala 43:32:@735.4]
  assign _GEN_21 = 7'h14 == _T_926 ? memory_20 : _GEN_20; // @[Mem.scala 43:32:@735.4]
  assign _GEN_22 = 7'h15 == _T_926 ? memory_21 : _GEN_21; // @[Mem.scala 43:32:@735.4]
  assign _GEN_23 = 7'h16 == _T_926 ? memory_22 : _GEN_22; // @[Mem.scala 43:32:@735.4]
  assign _GEN_24 = 7'h17 == _T_926 ? memory_23 : _GEN_23; // @[Mem.scala 43:32:@735.4]
  assign _GEN_25 = 7'h18 == _T_926 ? memory_24 : _GEN_24; // @[Mem.scala 43:32:@735.4]
  assign _GEN_26 = 7'h19 == _T_926 ? memory_25 : _GEN_25; // @[Mem.scala 43:32:@735.4]
  assign _GEN_27 = 7'h1a == _T_926 ? memory_26 : _GEN_26; // @[Mem.scala 43:32:@735.4]
  assign _GEN_28 = 7'h1b == _T_926 ? memory_27 : _GEN_27; // @[Mem.scala 43:32:@735.4]
  assign _GEN_29 = 7'h1c == _T_926 ? memory_28 : _GEN_28; // @[Mem.scala 43:32:@735.4]
  assign _GEN_30 = 7'h1d == _T_926 ? memory_29 : _GEN_29; // @[Mem.scala 43:32:@735.4]
  assign _GEN_31 = 7'h1e == _T_926 ? memory_30 : _GEN_30; // @[Mem.scala 43:32:@735.4]
  assign _GEN_32 = 7'h1f == _T_926 ? memory_31 : _GEN_31; // @[Mem.scala 43:32:@735.4]
  assign _GEN_33 = 7'h20 == _T_926 ? memory_32 : _GEN_32; // @[Mem.scala 43:32:@735.4]
  assign _GEN_34 = 7'h21 == _T_926 ? memory_33 : _GEN_33; // @[Mem.scala 43:32:@735.4]
  assign _GEN_35 = 7'h22 == _T_926 ? memory_34 : _GEN_34; // @[Mem.scala 43:32:@735.4]
  assign _GEN_36 = 7'h23 == _T_926 ? memory_35 : _GEN_35; // @[Mem.scala 43:32:@735.4]
  assign _GEN_37 = 7'h24 == _T_926 ? memory_36 : _GEN_36; // @[Mem.scala 43:32:@735.4]
  assign _GEN_38 = 7'h25 == _T_926 ? memory_37 : _GEN_37; // @[Mem.scala 43:32:@735.4]
  assign _GEN_39 = 7'h26 == _T_926 ? memory_38 : _GEN_38; // @[Mem.scala 43:32:@735.4]
  assign _GEN_40 = 7'h27 == _T_926 ? memory_39 : _GEN_39; // @[Mem.scala 43:32:@735.4]
  assign _GEN_41 = 7'h28 == _T_926 ? memory_40 : _GEN_40; // @[Mem.scala 43:32:@735.4]
  assign _GEN_42 = 7'h29 == _T_926 ? memory_41 : _GEN_41; // @[Mem.scala 43:32:@735.4]
  assign _GEN_43 = 7'h2a == _T_926 ? memory_42 : _GEN_42; // @[Mem.scala 43:32:@735.4]
  assign _GEN_44 = 7'h2b == _T_926 ? memory_43 : _GEN_43; // @[Mem.scala 43:32:@735.4]
  assign _GEN_45 = 7'h2c == _T_926 ? memory_44 : _GEN_44; // @[Mem.scala 43:32:@735.4]
  assign _GEN_46 = 7'h2d == _T_926 ? memory_45 : _GEN_45; // @[Mem.scala 43:32:@735.4]
  assign _GEN_47 = 7'h2e == _T_926 ? memory_46 : _GEN_46; // @[Mem.scala 43:32:@735.4]
  assign _GEN_48 = 7'h2f == _T_926 ? memory_47 : _GEN_47; // @[Mem.scala 43:32:@735.4]
  assign _GEN_49 = 7'h30 == _T_926 ? memory_48 : _GEN_48; // @[Mem.scala 43:32:@735.4]
  assign _GEN_50 = 7'h31 == _T_926 ? memory_49 : _GEN_49; // @[Mem.scala 43:32:@735.4]
  assign _GEN_51 = 7'h32 == _T_926 ? memory_50 : _GEN_50; // @[Mem.scala 43:32:@735.4]
  assign _GEN_52 = 7'h33 == _T_926 ? memory_51 : _GEN_51; // @[Mem.scala 43:32:@735.4]
  assign _GEN_53 = 7'h34 == _T_926 ? memory_52 : _GEN_52; // @[Mem.scala 43:32:@735.4]
  assign _GEN_54 = 7'h35 == _T_926 ? memory_53 : _GEN_53; // @[Mem.scala 43:32:@735.4]
  assign _GEN_55 = 7'h36 == _T_926 ? memory_54 : _GEN_54; // @[Mem.scala 43:32:@735.4]
  assign _GEN_56 = 7'h37 == _T_926 ? memory_55 : _GEN_55; // @[Mem.scala 43:32:@735.4]
  assign _GEN_57 = 7'h38 == _T_926 ? memory_56 : _GEN_56; // @[Mem.scala 43:32:@735.4]
  assign _GEN_58 = 7'h39 == _T_926 ? memory_57 : _GEN_57; // @[Mem.scala 43:32:@735.4]
  assign _GEN_59 = 7'h3a == _T_926 ? memory_58 : _GEN_58; // @[Mem.scala 43:32:@735.4]
  assign _GEN_60 = 7'h3b == _T_926 ? memory_59 : _GEN_59; // @[Mem.scala 43:32:@735.4]
  assign _GEN_61 = 7'h3c == _T_926 ? memory_60 : _GEN_60; // @[Mem.scala 43:32:@735.4]
  assign _GEN_62 = 7'h3d == _T_926 ? memory_61 : _GEN_61; // @[Mem.scala 43:32:@735.4]
  assign _GEN_63 = 7'h3e == _T_926 ? memory_62 : _GEN_62; // @[Mem.scala 43:32:@735.4]
  assign _GEN_64 = 7'h3f == _T_926 ? memory_63 : _GEN_63; // @[Mem.scala 43:32:@735.4]
  assign _GEN_65 = 7'h40 == _T_926 ? memory_64 : _GEN_64; // @[Mem.scala 43:32:@735.4]
  assign _GEN_66 = 7'h41 == _T_926 ? memory_65 : _GEN_65; // @[Mem.scala 43:32:@735.4]
  assign _GEN_67 = 7'h42 == _T_926 ? memory_66 : _GEN_66; // @[Mem.scala 43:32:@735.4]
  assign _GEN_68 = 7'h43 == _T_926 ? memory_67 : _GEN_67; // @[Mem.scala 43:32:@735.4]
  assign _GEN_69 = 7'h44 == _T_926 ? memory_68 : _GEN_68; // @[Mem.scala 43:32:@735.4]
  assign _GEN_70 = 7'h45 == _T_926 ? memory_69 : _GEN_69; // @[Mem.scala 43:32:@735.4]
  assign _GEN_71 = 7'h46 == _T_926 ? memory_70 : _GEN_70; // @[Mem.scala 43:32:@735.4]
  assign _GEN_72 = 7'h47 == _T_926 ? memory_71 : _GEN_71; // @[Mem.scala 43:32:@735.4]
  assign _GEN_73 = 7'h48 == _T_926 ? memory_72 : _GEN_72; // @[Mem.scala 43:32:@735.4]
  assign _GEN_74 = 7'h49 == _T_926 ? memory_73 : _GEN_73; // @[Mem.scala 43:32:@735.4]
  assign _GEN_75 = 7'h4a == _T_926 ? memory_74 : _GEN_74; // @[Mem.scala 43:32:@735.4]
  assign _GEN_76 = 7'h4b == _T_926 ? memory_75 : _GEN_75; // @[Mem.scala 43:32:@735.4]
  assign _GEN_77 = 7'h4c == _T_926 ? memory_76 : _GEN_76; // @[Mem.scala 43:32:@735.4]
  assign _GEN_78 = 7'h4d == _T_926 ? memory_77 : _GEN_77; // @[Mem.scala 43:32:@735.4]
  assign _GEN_79 = 7'h4e == _T_926 ? memory_78 : _GEN_78; // @[Mem.scala 43:32:@735.4]
  assign _GEN_80 = 7'h4f == _T_926 ? memory_79 : _GEN_79; // @[Mem.scala 43:32:@735.4]
  assign _GEN_81 = 7'h50 == _T_926 ? memory_80 : _GEN_80; // @[Mem.scala 43:32:@735.4]
  assign _GEN_82 = 7'h51 == _T_926 ? memory_81 : _GEN_81; // @[Mem.scala 43:32:@735.4]
  assign _GEN_83 = 7'h52 == _T_926 ? memory_82 : _GEN_82; // @[Mem.scala 43:32:@735.4]
  assign _GEN_84 = 7'h53 == _T_926 ? memory_83 : _GEN_83; // @[Mem.scala 43:32:@735.4]
  assign _GEN_85 = 7'h54 == _T_926 ? memory_84 : _GEN_84; // @[Mem.scala 43:32:@735.4]
  assign _GEN_86 = 7'h55 == _T_926 ? memory_85 : _GEN_85; // @[Mem.scala 43:32:@735.4]
  assign _GEN_87 = 7'h56 == _T_926 ? memory_86 : _GEN_86; // @[Mem.scala 43:32:@735.4]
  assign _GEN_88 = 7'h57 == _T_926 ? memory_87 : _GEN_87; // @[Mem.scala 43:32:@735.4]
  assign _GEN_89 = 7'h58 == _T_926 ? memory_88 : _GEN_88; // @[Mem.scala 43:32:@735.4]
  assign _GEN_90 = 7'h59 == _T_926 ? memory_89 : _GEN_89; // @[Mem.scala 43:32:@735.4]
  assign _GEN_91 = 7'h5a == _T_926 ? memory_90 : _GEN_90; // @[Mem.scala 43:32:@735.4]
  assign _GEN_92 = 7'h5b == _T_926 ? memory_91 : _GEN_91; // @[Mem.scala 43:32:@735.4]
  assign _GEN_93 = 7'h5c == _T_926 ? memory_92 : _GEN_92; // @[Mem.scala 43:32:@735.4]
  assign _GEN_94 = 7'h5d == _T_926 ? memory_93 : _GEN_93; // @[Mem.scala 43:32:@735.4]
  assign _GEN_95 = 7'h5e == _T_926 ? memory_94 : _GEN_94; // @[Mem.scala 43:32:@735.4]
  assign _GEN_96 = 7'h5f == _T_926 ? memory_95 : _GEN_95; // @[Mem.scala 43:32:@735.4]
  assign _GEN_97 = 7'h60 == _T_926 ? memory_96 : _GEN_96; // @[Mem.scala 43:32:@735.4]
  assign _GEN_98 = 7'h61 == _T_926 ? memory_97 : _GEN_97; // @[Mem.scala 43:32:@735.4]
  assign _GEN_99 = 7'h62 == _T_926 ? memory_98 : _GEN_98; // @[Mem.scala 43:32:@735.4]
  assign _GEN_100 = 7'h63 == _T_926 ? memory_99 : _GEN_99; // @[Mem.scala 43:32:@735.4]
  assign _GEN_101 = 7'h64 == _T_926 ? memory_100 : _GEN_100; // @[Mem.scala 43:32:@735.4]
  assign _GEN_102 = 7'h65 == _T_926 ? memory_101 : _GEN_101; // @[Mem.scala 43:32:@735.4]
  assign _GEN_103 = 7'h66 == _T_926 ? memory_102 : _GEN_102; // @[Mem.scala 43:32:@735.4]
  assign _GEN_104 = 7'h67 == _T_926 ? memory_103 : _GEN_103; // @[Mem.scala 43:32:@735.4]
  assign _GEN_105 = 7'h68 == _T_926 ? memory_104 : _GEN_104; // @[Mem.scala 43:32:@735.4]
  assign _GEN_106 = 7'h69 == _T_926 ? memory_105 : _GEN_105; // @[Mem.scala 43:32:@735.4]
  assign _GEN_107 = 7'h6a == _T_926 ? memory_106 : _GEN_106; // @[Mem.scala 43:32:@735.4]
  assign _GEN_108 = 7'h6b == _T_926 ? memory_107 : _GEN_107; // @[Mem.scala 43:32:@735.4]
  assign _GEN_109 = 7'h6c == _T_926 ? memory_108 : _GEN_108; // @[Mem.scala 43:32:@735.4]
  assign _GEN_110 = 7'h6d == _T_926 ? memory_109 : _GEN_109; // @[Mem.scala 43:32:@735.4]
  assign _GEN_111 = 7'h6e == _T_926 ? memory_110 : _GEN_110; // @[Mem.scala 43:32:@735.4]
  assign _GEN_112 = 7'h6f == _T_926 ? memory_111 : _GEN_111; // @[Mem.scala 43:32:@735.4]
  assign _GEN_113 = 7'h70 == _T_926 ? memory_112 : _GEN_112; // @[Mem.scala 43:32:@735.4]
  assign _GEN_114 = 7'h71 == _T_926 ? memory_113 : _GEN_113; // @[Mem.scala 43:32:@735.4]
  assign _GEN_115 = 7'h72 == _T_926 ? memory_114 : _GEN_114; // @[Mem.scala 43:32:@735.4]
  assign _GEN_116 = 7'h73 == _T_926 ? memory_115 : _GEN_115; // @[Mem.scala 43:32:@735.4]
  assign _GEN_117 = 7'h74 == _T_926 ? memory_116 : _GEN_116; // @[Mem.scala 43:32:@735.4]
  assign _GEN_118 = 7'h75 == _T_926 ? memory_117 : _GEN_117; // @[Mem.scala 43:32:@735.4]
  assign _GEN_119 = 7'h76 == _T_926 ? memory_118 : _GEN_118; // @[Mem.scala 43:32:@735.4]
  assign _GEN_120 = 7'h77 == _T_926 ? memory_119 : _GEN_119; // @[Mem.scala 43:32:@735.4]
  assign _GEN_121 = 7'h78 == _T_926 ? memory_120 : _GEN_120; // @[Mem.scala 43:32:@735.4]
  assign _GEN_122 = 7'h79 == _T_926 ? memory_121 : _GEN_121; // @[Mem.scala 43:32:@735.4]
  assign _GEN_123 = 7'h7a == _T_926 ? memory_122 : _GEN_122; // @[Mem.scala 43:32:@735.4]
  assign _GEN_124 = 7'h7b == _T_926 ? memory_123 : _GEN_123; // @[Mem.scala 43:32:@735.4]
  assign _GEN_125 = 7'h7c == _T_926 ? memory_124 : _GEN_124; // @[Mem.scala 43:32:@735.4]
  assign _GEN_126 = 7'h7d == _T_926 ? memory_125 : _GEN_125; // @[Mem.scala 43:32:@735.4]
  assign _GEN_127 = 7'h7e == _T_926 ? memory_126 : _GEN_126; // @[Mem.scala 43:32:@735.4]
  assign _T_930 = io_mem_addr == 32'h1; // @[Mem.scala 39:41:@737.4]
  assign _T_931 = io_mem_wen & _T_930; // @[Mem.scala 39:26:@738.4]
  assign _GEN_129 = _T_931 ? io_mem_wdata : memory_1; // @[Mem.scala 39:50:@739.4]
  assign _T_939 = io_mem_addr == 32'h2; // @[Mem.scala 39:41:@746.4]
  assign _T_940 = io_mem_wen & _T_939; // @[Mem.scala 39:26:@747.4]
  assign _GEN_258 = _T_940 ? io_mem_wdata : memory_2; // @[Mem.scala 39:50:@748.4]
  assign _T_948 = io_mem_addr == 32'h3; // @[Mem.scala 39:41:@755.4]
  assign _T_949 = io_mem_wen & _T_948; // @[Mem.scala 39:26:@756.4]
  assign _GEN_387 = _T_949 ? io_mem_wdata : memory_3; // @[Mem.scala 39:50:@757.4]
  assign _T_957 = io_mem_addr == 32'h4; // @[Mem.scala 39:41:@764.4]
  assign _T_958 = io_mem_wen & _T_957; // @[Mem.scala 39:26:@765.4]
  assign _GEN_516 = _T_958 ? io_mem_wdata : memory_4; // @[Mem.scala 39:50:@766.4]
  assign _T_966 = io_mem_addr == 32'h5; // @[Mem.scala 39:41:@773.4]
  assign _T_967 = io_mem_wen & _T_966; // @[Mem.scala 39:26:@774.4]
  assign _GEN_645 = _T_967 ? io_mem_wdata : memory_5; // @[Mem.scala 39:50:@775.4]
  assign _T_975 = io_mem_addr == 32'h6; // @[Mem.scala 39:41:@782.4]
  assign _T_976 = io_mem_wen & _T_975; // @[Mem.scala 39:26:@783.4]
  assign _GEN_774 = _T_976 ? io_mem_wdata : memory_6; // @[Mem.scala 39:50:@784.4]
  assign _T_984 = io_mem_addr == 32'h7; // @[Mem.scala 39:41:@791.4]
  assign _T_985 = io_mem_wen & _T_984; // @[Mem.scala 39:26:@792.4]
  assign _GEN_903 = _T_985 ? io_mem_wdata : memory_7; // @[Mem.scala 39:50:@793.4]
  assign _T_993 = io_mem_addr == 32'h8; // @[Mem.scala 39:41:@800.4]
  assign _T_994 = io_mem_wen & _T_993; // @[Mem.scala 39:26:@801.4]
  assign _GEN_1032 = _T_994 ? io_mem_wdata : memory_8; // @[Mem.scala 39:50:@802.4]
  assign _T_1002 = io_mem_addr == 32'h9; // @[Mem.scala 39:41:@809.4]
  assign _T_1003 = io_mem_wen & _T_1002; // @[Mem.scala 39:26:@810.4]
  assign _GEN_1161 = _T_1003 ? io_mem_wdata : memory_9; // @[Mem.scala 39:50:@811.4]
  assign _T_1011 = io_mem_addr == 32'ha; // @[Mem.scala 39:41:@818.4]
  assign _T_1012 = io_mem_wen & _T_1011; // @[Mem.scala 39:26:@819.4]
  assign _GEN_1290 = _T_1012 ? io_mem_wdata : memory_10; // @[Mem.scala 39:50:@820.4]
  assign _T_1020 = io_mem_addr == 32'hb; // @[Mem.scala 39:41:@827.4]
  assign _T_1021 = io_mem_wen & _T_1020; // @[Mem.scala 39:26:@828.4]
  assign _GEN_1419 = _T_1021 ? io_mem_wdata : memory_11; // @[Mem.scala 39:50:@829.4]
  assign _T_1029 = io_mem_addr == 32'hc; // @[Mem.scala 39:41:@836.4]
  assign _T_1030 = io_mem_wen & _T_1029; // @[Mem.scala 39:26:@837.4]
  assign _GEN_1548 = _T_1030 ? io_mem_wdata : memory_12; // @[Mem.scala 39:50:@838.4]
  assign _T_1038 = io_mem_addr == 32'hd; // @[Mem.scala 39:41:@845.4]
  assign _T_1039 = io_mem_wen & _T_1038; // @[Mem.scala 39:26:@846.4]
  assign _GEN_1677 = _T_1039 ? io_mem_wdata : memory_13; // @[Mem.scala 39:50:@847.4]
  assign _T_1047 = io_mem_addr == 32'he; // @[Mem.scala 39:41:@854.4]
  assign _T_1048 = io_mem_wen & _T_1047; // @[Mem.scala 39:26:@855.4]
  assign _GEN_1806 = _T_1048 ? io_mem_wdata : memory_14; // @[Mem.scala 39:50:@856.4]
  assign _T_1056 = io_mem_addr == 32'hf; // @[Mem.scala 39:41:@863.4]
  assign _T_1057 = io_mem_wen & _T_1056; // @[Mem.scala 39:26:@864.4]
  assign _GEN_1935 = _T_1057 ? io_mem_wdata : memory_15; // @[Mem.scala 39:50:@865.4]
  assign _T_1065 = io_mem_addr == 32'h10; // @[Mem.scala 39:41:@872.4]
  assign _T_1066 = io_mem_wen & _T_1065; // @[Mem.scala 39:26:@873.4]
  assign _GEN_2064 = _T_1066 ? io_mem_wdata : memory_16; // @[Mem.scala 39:50:@874.4]
  assign _T_1074 = io_mem_addr == 32'h11; // @[Mem.scala 39:41:@881.4]
  assign _T_1075 = io_mem_wen & _T_1074; // @[Mem.scala 39:26:@882.4]
  assign _GEN_2193 = _T_1075 ? io_mem_wdata : memory_17; // @[Mem.scala 39:50:@883.4]
  assign _T_1083 = io_mem_addr == 32'h12; // @[Mem.scala 39:41:@890.4]
  assign _T_1084 = io_mem_wen & _T_1083; // @[Mem.scala 39:26:@891.4]
  assign _GEN_2322 = _T_1084 ? io_mem_wdata : memory_18; // @[Mem.scala 39:50:@892.4]
  assign _T_1092 = io_mem_addr == 32'h13; // @[Mem.scala 39:41:@899.4]
  assign _T_1093 = io_mem_wen & _T_1092; // @[Mem.scala 39:26:@900.4]
  assign _GEN_2451 = _T_1093 ? io_mem_wdata : memory_19; // @[Mem.scala 39:50:@901.4]
  assign _T_1101 = io_mem_addr == 32'h14; // @[Mem.scala 39:41:@908.4]
  assign _T_1102 = io_mem_wen & _T_1101; // @[Mem.scala 39:26:@909.4]
  assign _GEN_2580 = _T_1102 ? io_mem_wdata : memory_20; // @[Mem.scala 39:50:@910.4]
  assign _T_1110 = io_mem_addr == 32'h15; // @[Mem.scala 39:41:@917.4]
  assign _T_1111 = io_mem_wen & _T_1110; // @[Mem.scala 39:26:@918.4]
  assign _GEN_2709 = _T_1111 ? io_mem_wdata : memory_21; // @[Mem.scala 39:50:@919.4]
  assign _T_1119 = io_mem_addr == 32'h16; // @[Mem.scala 39:41:@926.4]
  assign _T_1120 = io_mem_wen & _T_1119; // @[Mem.scala 39:26:@927.4]
  assign _GEN_2838 = _T_1120 ? io_mem_wdata : memory_22; // @[Mem.scala 39:50:@928.4]
  assign _T_1128 = io_mem_addr == 32'h17; // @[Mem.scala 39:41:@935.4]
  assign _T_1129 = io_mem_wen & _T_1128; // @[Mem.scala 39:26:@936.4]
  assign _GEN_2967 = _T_1129 ? io_mem_wdata : memory_23; // @[Mem.scala 39:50:@937.4]
  assign _T_1137 = io_mem_addr == 32'h18; // @[Mem.scala 39:41:@944.4]
  assign _T_1138 = io_mem_wen & _T_1137; // @[Mem.scala 39:26:@945.4]
  assign _GEN_3096 = _T_1138 ? io_mem_wdata : memory_24; // @[Mem.scala 39:50:@946.4]
  assign _T_1146 = io_mem_addr == 32'h19; // @[Mem.scala 39:41:@953.4]
  assign _T_1147 = io_mem_wen & _T_1146; // @[Mem.scala 39:26:@954.4]
  assign _GEN_3225 = _T_1147 ? io_mem_wdata : memory_25; // @[Mem.scala 39:50:@955.4]
  assign _T_1155 = io_mem_addr == 32'h1a; // @[Mem.scala 39:41:@962.4]
  assign _T_1156 = io_mem_wen & _T_1155; // @[Mem.scala 39:26:@963.4]
  assign _GEN_3354 = _T_1156 ? io_mem_wdata : memory_26; // @[Mem.scala 39:50:@964.4]
  assign _T_1164 = io_mem_addr == 32'h1b; // @[Mem.scala 39:41:@971.4]
  assign _T_1165 = io_mem_wen & _T_1164; // @[Mem.scala 39:26:@972.4]
  assign _GEN_3483 = _T_1165 ? io_mem_wdata : memory_27; // @[Mem.scala 39:50:@973.4]
  assign _T_1173 = io_mem_addr == 32'h1c; // @[Mem.scala 39:41:@980.4]
  assign _T_1174 = io_mem_wen & _T_1173; // @[Mem.scala 39:26:@981.4]
  assign _GEN_3612 = _T_1174 ? io_mem_wdata : memory_28; // @[Mem.scala 39:50:@982.4]
  assign _T_1182 = io_mem_addr == 32'h1d; // @[Mem.scala 39:41:@989.4]
  assign _T_1183 = io_mem_wen & _T_1182; // @[Mem.scala 39:26:@990.4]
  assign _GEN_3741 = _T_1183 ? io_mem_wdata : memory_29; // @[Mem.scala 39:50:@991.4]
  assign _T_1191 = io_mem_addr == 32'h1e; // @[Mem.scala 39:41:@998.4]
  assign _T_1192 = io_mem_wen & _T_1191; // @[Mem.scala 39:26:@999.4]
  assign _GEN_3870 = _T_1192 ? io_mem_wdata : memory_30; // @[Mem.scala 39:50:@1000.4]
  assign _T_1200 = io_mem_addr == 32'h1f; // @[Mem.scala 39:41:@1007.4]
  assign _T_1201 = io_mem_wen & _T_1200; // @[Mem.scala 39:26:@1008.4]
  assign _GEN_3999 = _T_1201 ? io_mem_wdata : memory_31; // @[Mem.scala 39:50:@1009.4]
  assign _T_1209 = io_mem_addr == 32'h20; // @[Mem.scala 39:41:@1016.4]
  assign _T_1210 = io_mem_wen & _T_1209; // @[Mem.scala 39:26:@1017.4]
  assign _GEN_4128 = _T_1210 ? io_mem_wdata : memory_32; // @[Mem.scala 39:50:@1018.4]
  assign _T_1218 = io_mem_addr == 32'h21; // @[Mem.scala 39:41:@1025.4]
  assign _T_1219 = io_mem_wen & _T_1218; // @[Mem.scala 39:26:@1026.4]
  assign _GEN_4257 = _T_1219 ? io_mem_wdata : memory_33; // @[Mem.scala 39:50:@1027.4]
  assign _T_1227 = io_mem_addr == 32'h22; // @[Mem.scala 39:41:@1034.4]
  assign _T_1228 = io_mem_wen & _T_1227; // @[Mem.scala 39:26:@1035.4]
  assign _GEN_4386 = _T_1228 ? io_mem_wdata : memory_34; // @[Mem.scala 39:50:@1036.4]
  assign _T_1236 = io_mem_addr == 32'h23; // @[Mem.scala 39:41:@1043.4]
  assign _T_1237 = io_mem_wen & _T_1236; // @[Mem.scala 39:26:@1044.4]
  assign _GEN_4515 = _T_1237 ? io_mem_wdata : memory_35; // @[Mem.scala 39:50:@1045.4]
  assign _T_1245 = io_mem_addr == 32'h24; // @[Mem.scala 39:41:@1052.4]
  assign _T_1246 = io_mem_wen & _T_1245; // @[Mem.scala 39:26:@1053.4]
  assign _GEN_4644 = _T_1246 ? io_mem_wdata : memory_36; // @[Mem.scala 39:50:@1054.4]
  assign _T_1254 = io_mem_addr == 32'h25; // @[Mem.scala 39:41:@1061.4]
  assign _T_1255 = io_mem_wen & _T_1254; // @[Mem.scala 39:26:@1062.4]
  assign _GEN_4773 = _T_1255 ? io_mem_wdata : memory_37; // @[Mem.scala 39:50:@1063.4]
  assign _T_1263 = io_mem_addr == 32'h26; // @[Mem.scala 39:41:@1070.4]
  assign _T_1264 = io_mem_wen & _T_1263; // @[Mem.scala 39:26:@1071.4]
  assign _GEN_4902 = _T_1264 ? io_mem_wdata : memory_38; // @[Mem.scala 39:50:@1072.4]
  assign _T_1272 = io_mem_addr == 32'h27; // @[Mem.scala 39:41:@1079.4]
  assign _T_1273 = io_mem_wen & _T_1272; // @[Mem.scala 39:26:@1080.4]
  assign _GEN_5031 = _T_1273 ? io_mem_wdata : memory_39; // @[Mem.scala 39:50:@1081.4]
  assign _T_1281 = io_mem_addr == 32'h28; // @[Mem.scala 39:41:@1088.4]
  assign _T_1282 = io_mem_wen & _T_1281; // @[Mem.scala 39:26:@1089.4]
  assign _GEN_5160 = _T_1282 ? io_mem_wdata : memory_40; // @[Mem.scala 39:50:@1090.4]
  assign _T_1290 = io_mem_addr == 32'h29; // @[Mem.scala 39:41:@1097.4]
  assign _T_1291 = io_mem_wen & _T_1290; // @[Mem.scala 39:26:@1098.4]
  assign _GEN_5289 = _T_1291 ? io_mem_wdata : memory_41; // @[Mem.scala 39:50:@1099.4]
  assign _T_1299 = io_mem_addr == 32'h2a; // @[Mem.scala 39:41:@1106.4]
  assign _T_1300 = io_mem_wen & _T_1299; // @[Mem.scala 39:26:@1107.4]
  assign _GEN_5418 = _T_1300 ? io_mem_wdata : memory_42; // @[Mem.scala 39:50:@1108.4]
  assign _T_1308 = io_mem_addr == 32'h2b; // @[Mem.scala 39:41:@1115.4]
  assign _T_1309 = io_mem_wen & _T_1308; // @[Mem.scala 39:26:@1116.4]
  assign _GEN_5547 = _T_1309 ? io_mem_wdata : memory_43; // @[Mem.scala 39:50:@1117.4]
  assign _T_1317 = io_mem_addr == 32'h2c; // @[Mem.scala 39:41:@1124.4]
  assign _T_1318 = io_mem_wen & _T_1317; // @[Mem.scala 39:26:@1125.4]
  assign _GEN_5676 = _T_1318 ? io_mem_wdata : memory_44; // @[Mem.scala 39:50:@1126.4]
  assign _T_1326 = io_mem_addr == 32'h2d; // @[Mem.scala 39:41:@1133.4]
  assign _T_1327 = io_mem_wen & _T_1326; // @[Mem.scala 39:26:@1134.4]
  assign _GEN_5805 = _T_1327 ? io_mem_wdata : memory_45; // @[Mem.scala 39:50:@1135.4]
  assign _T_1335 = io_mem_addr == 32'h2e; // @[Mem.scala 39:41:@1142.4]
  assign _T_1336 = io_mem_wen & _T_1335; // @[Mem.scala 39:26:@1143.4]
  assign _GEN_5934 = _T_1336 ? io_mem_wdata : memory_46; // @[Mem.scala 39:50:@1144.4]
  assign _T_1344 = io_mem_addr == 32'h2f; // @[Mem.scala 39:41:@1151.4]
  assign _T_1345 = io_mem_wen & _T_1344; // @[Mem.scala 39:26:@1152.4]
  assign _GEN_6063 = _T_1345 ? io_mem_wdata : memory_47; // @[Mem.scala 39:50:@1153.4]
  assign _T_1353 = io_mem_addr == 32'h30; // @[Mem.scala 39:41:@1160.4]
  assign _T_1354 = io_mem_wen & _T_1353; // @[Mem.scala 39:26:@1161.4]
  assign _GEN_6192 = _T_1354 ? io_mem_wdata : memory_48; // @[Mem.scala 39:50:@1162.4]
  assign _T_1362 = io_mem_addr == 32'h31; // @[Mem.scala 39:41:@1169.4]
  assign _T_1363 = io_mem_wen & _T_1362; // @[Mem.scala 39:26:@1170.4]
  assign _GEN_6321 = _T_1363 ? io_mem_wdata : memory_49; // @[Mem.scala 39:50:@1171.4]
  assign _T_1371 = io_mem_addr == 32'h32; // @[Mem.scala 39:41:@1178.4]
  assign _T_1372 = io_mem_wen & _T_1371; // @[Mem.scala 39:26:@1179.4]
  assign _GEN_6450 = _T_1372 ? io_mem_wdata : memory_50; // @[Mem.scala 39:50:@1180.4]
  assign _T_1380 = io_mem_addr == 32'h33; // @[Mem.scala 39:41:@1187.4]
  assign _T_1381 = io_mem_wen & _T_1380; // @[Mem.scala 39:26:@1188.4]
  assign _GEN_6579 = _T_1381 ? io_mem_wdata : memory_51; // @[Mem.scala 39:50:@1189.4]
  assign _T_1389 = io_mem_addr == 32'h34; // @[Mem.scala 39:41:@1196.4]
  assign _T_1390 = io_mem_wen & _T_1389; // @[Mem.scala 39:26:@1197.4]
  assign _GEN_6708 = _T_1390 ? io_mem_wdata : memory_52; // @[Mem.scala 39:50:@1198.4]
  assign _T_1398 = io_mem_addr == 32'h35; // @[Mem.scala 39:41:@1205.4]
  assign _T_1399 = io_mem_wen & _T_1398; // @[Mem.scala 39:26:@1206.4]
  assign _GEN_6837 = _T_1399 ? io_mem_wdata : memory_53; // @[Mem.scala 39:50:@1207.4]
  assign _T_1407 = io_mem_addr == 32'h36; // @[Mem.scala 39:41:@1214.4]
  assign _T_1408 = io_mem_wen & _T_1407; // @[Mem.scala 39:26:@1215.4]
  assign _GEN_6966 = _T_1408 ? io_mem_wdata : memory_54; // @[Mem.scala 39:50:@1216.4]
  assign _T_1416 = io_mem_addr == 32'h37; // @[Mem.scala 39:41:@1223.4]
  assign _T_1417 = io_mem_wen & _T_1416; // @[Mem.scala 39:26:@1224.4]
  assign _GEN_7095 = _T_1417 ? io_mem_wdata : memory_55; // @[Mem.scala 39:50:@1225.4]
  assign _T_1425 = io_mem_addr == 32'h38; // @[Mem.scala 39:41:@1232.4]
  assign _T_1426 = io_mem_wen & _T_1425; // @[Mem.scala 39:26:@1233.4]
  assign _GEN_7224 = _T_1426 ? io_mem_wdata : memory_56; // @[Mem.scala 39:50:@1234.4]
  assign _T_1434 = io_mem_addr == 32'h39; // @[Mem.scala 39:41:@1241.4]
  assign _T_1435 = io_mem_wen & _T_1434; // @[Mem.scala 39:26:@1242.4]
  assign _GEN_7353 = _T_1435 ? io_mem_wdata : memory_57; // @[Mem.scala 39:50:@1243.4]
  assign _T_1443 = io_mem_addr == 32'h3a; // @[Mem.scala 39:41:@1250.4]
  assign _T_1444 = io_mem_wen & _T_1443; // @[Mem.scala 39:26:@1251.4]
  assign _GEN_7482 = _T_1444 ? io_mem_wdata : memory_58; // @[Mem.scala 39:50:@1252.4]
  assign _T_1452 = io_mem_addr == 32'h3b; // @[Mem.scala 39:41:@1259.4]
  assign _T_1453 = io_mem_wen & _T_1452; // @[Mem.scala 39:26:@1260.4]
  assign _GEN_7611 = _T_1453 ? io_mem_wdata : memory_59; // @[Mem.scala 39:50:@1261.4]
  assign _T_1461 = io_mem_addr == 32'h3c; // @[Mem.scala 39:41:@1268.4]
  assign _T_1462 = io_mem_wen & _T_1461; // @[Mem.scala 39:26:@1269.4]
  assign _GEN_7740 = _T_1462 ? io_mem_wdata : memory_60; // @[Mem.scala 39:50:@1270.4]
  assign _T_1470 = io_mem_addr == 32'h3d; // @[Mem.scala 39:41:@1277.4]
  assign _T_1471 = io_mem_wen & _T_1470; // @[Mem.scala 39:26:@1278.4]
  assign _GEN_7869 = _T_1471 ? io_mem_wdata : memory_61; // @[Mem.scala 39:50:@1279.4]
  assign _T_1479 = io_mem_addr == 32'h3e; // @[Mem.scala 39:41:@1286.4]
  assign _T_1480 = io_mem_wen & _T_1479; // @[Mem.scala 39:26:@1287.4]
  assign _GEN_7998 = _T_1480 ? io_mem_wdata : memory_62; // @[Mem.scala 39:50:@1288.4]
  assign _T_1488 = io_mem_addr == 32'h3f; // @[Mem.scala 39:41:@1295.4]
  assign _T_1489 = io_mem_wen & _T_1488; // @[Mem.scala 39:26:@1296.4]
  assign _GEN_8127 = _T_1489 ? io_mem_wdata : memory_63; // @[Mem.scala 39:50:@1297.4]
  assign _T_1497 = io_mem_addr == 32'h40; // @[Mem.scala 39:41:@1304.4]
  assign _T_1498 = io_mem_wen & _T_1497; // @[Mem.scala 39:26:@1305.4]
  assign _GEN_8256 = _T_1498 ? io_mem_wdata : memory_64; // @[Mem.scala 39:50:@1306.4]
  assign _T_1506 = io_mem_addr == 32'h41; // @[Mem.scala 39:41:@1313.4]
  assign _T_1507 = io_mem_wen & _T_1506; // @[Mem.scala 39:26:@1314.4]
  assign _GEN_8385 = _T_1507 ? io_mem_wdata : memory_65; // @[Mem.scala 39:50:@1315.4]
  assign _T_1515 = io_mem_addr == 32'h42; // @[Mem.scala 39:41:@1322.4]
  assign _T_1516 = io_mem_wen & _T_1515; // @[Mem.scala 39:26:@1323.4]
  assign _GEN_8514 = _T_1516 ? io_mem_wdata : memory_66; // @[Mem.scala 39:50:@1324.4]
  assign _T_1524 = io_mem_addr == 32'h43; // @[Mem.scala 39:41:@1331.4]
  assign _T_1525 = io_mem_wen & _T_1524; // @[Mem.scala 39:26:@1332.4]
  assign _GEN_8643 = _T_1525 ? io_mem_wdata : memory_67; // @[Mem.scala 39:50:@1333.4]
  assign _T_1533 = io_mem_addr == 32'h44; // @[Mem.scala 39:41:@1340.4]
  assign _T_1534 = io_mem_wen & _T_1533; // @[Mem.scala 39:26:@1341.4]
  assign _GEN_8772 = _T_1534 ? io_mem_wdata : memory_68; // @[Mem.scala 39:50:@1342.4]
  assign _T_1542 = io_mem_addr == 32'h45; // @[Mem.scala 39:41:@1349.4]
  assign _T_1543 = io_mem_wen & _T_1542; // @[Mem.scala 39:26:@1350.4]
  assign _GEN_8901 = _T_1543 ? io_mem_wdata : memory_69; // @[Mem.scala 39:50:@1351.4]
  assign _T_1551 = io_mem_addr == 32'h46; // @[Mem.scala 39:41:@1358.4]
  assign _T_1552 = io_mem_wen & _T_1551; // @[Mem.scala 39:26:@1359.4]
  assign _GEN_9030 = _T_1552 ? io_mem_wdata : memory_70; // @[Mem.scala 39:50:@1360.4]
  assign _T_1560 = io_mem_addr == 32'h47; // @[Mem.scala 39:41:@1367.4]
  assign _T_1561 = io_mem_wen & _T_1560; // @[Mem.scala 39:26:@1368.4]
  assign _GEN_9159 = _T_1561 ? io_mem_wdata : memory_71; // @[Mem.scala 39:50:@1369.4]
  assign _T_1569 = io_mem_addr == 32'h48; // @[Mem.scala 39:41:@1376.4]
  assign _T_1570 = io_mem_wen & _T_1569; // @[Mem.scala 39:26:@1377.4]
  assign _GEN_9288 = _T_1570 ? io_mem_wdata : memory_72; // @[Mem.scala 39:50:@1378.4]
  assign _T_1578 = io_mem_addr == 32'h49; // @[Mem.scala 39:41:@1385.4]
  assign _T_1579 = io_mem_wen & _T_1578; // @[Mem.scala 39:26:@1386.4]
  assign _GEN_9417 = _T_1579 ? io_mem_wdata : memory_73; // @[Mem.scala 39:50:@1387.4]
  assign _T_1587 = io_mem_addr == 32'h4a; // @[Mem.scala 39:41:@1394.4]
  assign _T_1588 = io_mem_wen & _T_1587; // @[Mem.scala 39:26:@1395.4]
  assign _GEN_9546 = _T_1588 ? io_mem_wdata : memory_74; // @[Mem.scala 39:50:@1396.4]
  assign _T_1596 = io_mem_addr == 32'h4b; // @[Mem.scala 39:41:@1403.4]
  assign _T_1597 = io_mem_wen & _T_1596; // @[Mem.scala 39:26:@1404.4]
  assign _GEN_9675 = _T_1597 ? io_mem_wdata : memory_75; // @[Mem.scala 39:50:@1405.4]
  assign _T_1605 = io_mem_addr == 32'h4c; // @[Mem.scala 39:41:@1412.4]
  assign _T_1606 = io_mem_wen & _T_1605; // @[Mem.scala 39:26:@1413.4]
  assign _GEN_9804 = _T_1606 ? io_mem_wdata : memory_76; // @[Mem.scala 39:50:@1414.4]
  assign _T_1614 = io_mem_addr == 32'h4d; // @[Mem.scala 39:41:@1421.4]
  assign _T_1615 = io_mem_wen & _T_1614; // @[Mem.scala 39:26:@1422.4]
  assign _GEN_9933 = _T_1615 ? io_mem_wdata : memory_77; // @[Mem.scala 39:50:@1423.4]
  assign _T_1623 = io_mem_addr == 32'h4e; // @[Mem.scala 39:41:@1430.4]
  assign _T_1624 = io_mem_wen & _T_1623; // @[Mem.scala 39:26:@1431.4]
  assign _GEN_10062 = _T_1624 ? io_mem_wdata : memory_78; // @[Mem.scala 39:50:@1432.4]
  assign _T_1632 = io_mem_addr == 32'h4f; // @[Mem.scala 39:41:@1439.4]
  assign _T_1633 = io_mem_wen & _T_1632; // @[Mem.scala 39:26:@1440.4]
  assign _GEN_10191 = _T_1633 ? io_mem_wdata : memory_79; // @[Mem.scala 39:50:@1441.4]
  assign _T_1641 = io_mem_addr == 32'h50; // @[Mem.scala 39:41:@1448.4]
  assign _T_1642 = io_mem_wen & _T_1641; // @[Mem.scala 39:26:@1449.4]
  assign _GEN_10320 = _T_1642 ? io_mem_wdata : memory_80; // @[Mem.scala 39:50:@1450.4]
  assign _T_1650 = io_mem_addr == 32'h51; // @[Mem.scala 39:41:@1457.4]
  assign _T_1651 = io_mem_wen & _T_1650; // @[Mem.scala 39:26:@1458.4]
  assign _GEN_10449 = _T_1651 ? io_mem_wdata : memory_81; // @[Mem.scala 39:50:@1459.4]
  assign _T_1659 = io_mem_addr == 32'h52; // @[Mem.scala 39:41:@1466.4]
  assign _T_1660 = io_mem_wen & _T_1659; // @[Mem.scala 39:26:@1467.4]
  assign _GEN_10578 = _T_1660 ? io_mem_wdata : memory_82; // @[Mem.scala 39:50:@1468.4]
  assign _T_1668 = io_mem_addr == 32'h53; // @[Mem.scala 39:41:@1475.4]
  assign _T_1669 = io_mem_wen & _T_1668; // @[Mem.scala 39:26:@1476.4]
  assign _GEN_10707 = _T_1669 ? io_mem_wdata : memory_83; // @[Mem.scala 39:50:@1477.4]
  assign _T_1677 = io_mem_addr == 32'h54; // @[Mem.scala 39:41:@1484.4]
  assign _T_1678 = io_mem_wen & _T_1677; // @[Mem.scala 39:26:@1485.4]
  assign _GEN_10836 = _T_1678 ? io_mem_wdata : memory_84; // @[Mem.scala 39:50:@1486.4]
  assign _T_1686 = io_mem_addr == 32'h55; // @[Mem.scala 39:41:@1493.4]
  assign _T_1687 = io_mem_wen & _T_1686; // @[Mem.scala 39:26:@1494.4]
  assign _GEN_10965 = _T_1687 ? io_mem_wdata : memory_85; // @[Mem.scala 39:50:@1495.4]
  assign _T_1695 = io_mem_addr == 32'h56; // @[Mem.scala 39:41:@1502.4]
  assign _T_1696 = io_mem_wen & _T_1695; // @[Mem.scala 39:26:@1503.4]
  assign _GEN_11094 = _T_1696 ? io_mem_wdata : memory_86; // @[Mem.scala 39:50:@1504.4]
  assign _T_1704 = io_mem_addr == 32'h57; // @[Mem.scala 39:41:@1511.4]
  assign _T_1705 = io_mem_wen & _T_1704; // @[Mem.scala 39:26:@1512.4]
  assign _GEN_11223 = _T_1705 ? io_mem_wdata : memory_87; // @[Mem.scala 39:50:@1513.4]
  assign _T_1713 = io_mem_addr == 32'h58; // @[Mem.scala 39:41:@1520.4]
  assign _T_1714 = io_mem_wen & _T_1713; // @[Mem.scala 39:26:@1521.4]
  assign _GEN_11352 = _T_1714 ? io_mem_wdata : memory_88; // @[Mem.scala 39:50:@1522.4]
  assign _T_1722 = io_mem_addr == 32'h59; // @[Mem.scala 39:41:@1529.4]
  assign _T_1723 = io_mem_wen & _T_1722; // @[Mem.scala 39:26:@1530.4]
  assign _GEN_11481 = _T_1723 ? io_mem_wdata : memory_89; // @[Mem.scala 39:50:@1531.4]
  assign _T_1731 = io_mem_addr == 32'h5a; // @[Mem.scala 39:41:@1538.4]
  assign _T_1732 = io_mem_wen & _T_1731; // @[Mem.scala 39:26:@1539.4]
  assign _GEN_11610 = _T_1732 ? io_mem_wdata : memory_90; // @[Mem.scala 39:50:@1540.4]
  assign _T_1740 = io_mem_addr == 32'h5b; // @[Mem.scala 39:41:@1547.4]
  assign _T_1741 = io_mem_wen & _T_1740; // @[Mem.scala 39:26:@1548.4]
  assign _GEN_11739 = _T_1741 ? io_mem_wdata : memory_91; // @[Mem.scala 39:50:@1549.4]
  assign _T_1749 = io_mem_addr == 32'h5c; // @[Mem.scala 39:41:@1556.4]
  assign _T_1750 = io_mem_wen & _T_1749; // @[Mem.scala 39:26:@1557.4]
  assign _GEN_11868 = _T_1750 ? io_mem_wdata : memory_92; // @[Mem.scala 39:50:@1558.4]
  assign _T_1758 = io_mem_addr == 32'h5d; // @[Mem.scala 39:41:@1565.4]
  assign _T_1759 = io_mem_wen & _T_1758; // @[Mem.scala 39:26:@1566.4]
  assign _GEN_11997 = _T_1759 ? io_mem_wdata : memory_93; // @[Mem.scala 39:50:@1567.4]
  assign _T_1767 = io_mem_addr == 32'h5e; // @[Mem.scala 39:41:@1574.4]
  assign _T_1768 = io_mem_wen & _T_1767; // @[Mem.scala 39:26:@1575.4]
  assign _GEN_12126 = _T_1768 ? io_mem_wdata : memory_94; // @[Mem.scala 39:50:@1576.4]
  assign _T_1776 = io_mem_addr == 32'h5f; // @[Mem.scala 39:41:@1583.4]
  assign _T_1777 = io_mem_wen & _T_1776; // @[Mem.scala 39:26:@1584.4]
  assign _GEN_12255 = _T_1777 ? io_mem_wdata : memory_95; // @[Mem.scala 39:50:@1585.4]
  assign _T_1785 = io_mem_addr == 32'h60; // @[Mem.scala 39:41:@1592.4]
  assign _T_1786 = io_mem_wen & _T_1785; // @[Mem.scala 39:26:@1593.4]
  assign _GEN_12384 = _T_1786 ? io_mem_wdata : memory_96; // @[Mem.scala 39:50:@1594.4]
  assign _T_1794 = io_mem_addr == 32'h61; // @[Mem.scala 39:41:@1601.4]
  assign _T_1795 = io_mem_wen & _T_1794; // @[Mem.scala 39:26:@1602.4]
  assign _GEN_12513 = _T_1795 ? io_mem_wdata : memory_97; // @[Mem.scala 39:50:@1603.4]
  assign _T_1803 = io_mem_addr == 32'h62; // @[Mem.scala 39:41:@1610.4]
  assign _T_1804 = io_mem_wen & _T_1803; // @[Mem.scala 39:26:@1611.4]
  assign _GEN_12642 = _T_1804 ? io_mem_wdata : memory_98; // @[Mem.scala 39:50:@1612.4]
  assign _T_1812 = io_mem_addr == 32'h63; // @[Mem.scala 39:41:@1619.4]
  assign _T_1813 = io_mem_wen & _T_1812; // @[Mem.scala 39:26:@1620.4]
  assign _GEN_12771 = _T_1813 ? io_mem_wdata : memory_99; // @[Mem.scala 39:50:@1621.4]
  assign _T_1821 = io_mem_addr == 32'h64; // @[Mem.scala 39:41:@1628.4]
  assign _T_1822 = io_mem_wen & _T_1821; // @[Mem.scala 39:26:@1629.4]
  assign _GEN_12900 = _T_1822 ? io_mem_wdata : memory_100; // @[Mem.scala 39:50:@1630.4]
  assign _T_1830 = io_mem_addr == 32'h65; // @[Mem.scala 39:41:@1637.4]
  assign _T_1831 = io_mem_wen & _T_1830; // @[Mem.scala 39:26:@1638.4]
  assign _GEN_13029 = _T_1831 ? io_mem_wdata : memory_101; // @[Mem.scala 39:50:@1639.4]
  assign _T_1839 = io_mem_addr == 32'h66; // @[Mem.scala 39:41:@1646.4]
  assign _T_1840 = io_mem_wen & _T_1839; // @[Mem.scala 39:26:@1647.4]
  assign _GEN_13158 = _T_1840 ? io_mem_wdata : memory_102; // @[Mem.scala 39:50:@1648.4]
  assign _T_1848 = io_mem_addr == 32'h67; // @[Mem.scala 39:41:@1655.4]
  assign _T_1849 = io_mem_wen & _T_1848; // @[Mem.scala 39:26:@1656.4]
  assign _GEN_13287 = _T_1849 ? io_mem_wdata : memory_103; // @[Mem.scala 39:50:@1657.4]
  assign _T_1857 = io_mem_addr == 32'h68; // @[Mem.scala 39:41:@1664.4]
  assign _T_1858 = io_mem_wen & _T_1857; // @[Mem.scala 39:26:@1665.4]
  assign _GEN_13416 = _T_1858 ? io_mem_wdata : memory_104; // @[Mem.scala 39:50:@1666.4]
  assign _T_1866 = io_mem_addr == 32'h69; // @[Mem.scala 39:41:@1673.4]
  assign _T_1867 = io_mem_wen & _T_1866; // @[Mem.scala 39:26:@1674.4]
  assign _GEN_13545 = _T_1867 ? io_mem_wdata : memory_105; // @[Mem.scala 39:50:@1675.4]
  assign _T_1875 = io_mem_addr == 32'h6a; // @[Mem.scala 39:41:@1682.4]
  assign _T_1876 = io_mem_wen & _T_1875; // @[Mem.scala 39:26:@1683.4]
  assign _GEN_13674 = _T_1876 ? io_mem_wdata : memory_106; // @[Mem.scala 39:50:@1684.4]
  assign _T_1884 = io_mem_addr == 32'h6b; // @[Mem.scala 39:41:@1691.4]
  assign _T_1885 = io_mem_wen & _T_1884; // @[Mem.scala 39:26:@1692.4]
  assign _GEN_13803 = _T_1885 ? io_mem_wdata : memory_107; // @[Mem.scala 39:50:@1693.4]
  assign _T_1893 = io_mem_addr == 32'h6c; // @[Mem.scala 39:41:@1700.4]
  assign _T_1894 = io_mem_wen & _T_1893; // @[Mem.scala 39:26:@1701.4]
  assign _GEN_13932 = _T_1894 ? io_mem_wdata : memory_108; // @[Mem.scala 39:50:@1702.4]
  assign _T_1902 = io_mem_addr == 32'h6d; // @[Mem.scala 39:41:@1709.4]
  assign _T_1903 = io_mem_wen & _T_1902; // @[Mem.scala 39:26:@1710.4]
  assign _GEN_14061 = _T_1903 ? io_mem_wdata : memory_109; // @[Mem.scala 39:50:@1711.4]
  assign _T_1911 = io_mem_addr == 32'h6e; // @[Mem.scala 39:41:@1718.4]
  assign _T_1912 = io_mem_wen & _T_1911; // @[Mem.scala 39:26:@1719.4]
  assign _GEN_14190 = _T_1912 ? io_mem_wdata : memory_110; // @[Mem.scala 39:50:@1720.4]
  assign _T_1920 = io_mem_addr == 32'h6f; // @[Mem.scala 39:41:@1727.4]
  assign _T_1921 = io_mem_wen & _T_1920; // @[Mem.scala 39:26:@1728.4]
  assign _GEN_14319 = _T_1921 ? io_mem_wdata : memory_111; // @[Mem.scala 39:50:@1729.4]
  assign _T_1929 = io_mem_addr == 32'h70; // @[Mem.scala 39:41:@1736.4]
  assign _T_1930 = io_mem_wen & _T_1929; // @[Mem.scala 39:26:@1737.4]
  assign _GEN_14448 = _T_1930 ? io_mem_wdata : memory_112; // @[Mem.scala 39:50:@1738.4]
  assign _T_1938 = io_mem_addr == 32'h71; // @[Mem.scala 39:41:@1745.4]
  assign _T_1939 = io_mem_wen & _T_1938; // @[Mem.scala 39:26:@1746.4]
  assign _GEN_14577 = _T_1939 ? io_mem_wdata : memory_113; // @[Mem.scala 39:50:@1747.4]
  assign _T_1947 = io_mem_addr == 32'h72; // @[Mem.scala 39:41:@1754.4]
  assign _T_1948 = io_mem_wen & _T_1947; // @[Mem.scala 39:26:@1755.4]
  assign _GEN_14706 = _T_1948 ? io_mem_wdata : memory_114; // @[Mem.scala 39:50:@1756.4]
  assign _T_1956 = io_mem_addr == 32'h73; // @[Mem.scala 39:41:@1763.4]
  assign _T_1957 = io_mem_wen & _T_1956; // @[Mem.scala 39:26:@1764.4]
  assign _GEN_14835 = _T_1957 ? io_mem_wdata : memory_115; // @[Mem.scala 39:50:@1765.4]
  assign _T_1965 = io_mem_addr == 32'h74; // @[Mem.scala 39:41:@1772.4]
  assign _T_1966 = io_mem_wen & _T_1965; // @[Mem.scala 39:26:@1773.4]
  assign _GEN_14964 = _T_1966 ? io_mem_wdata : memory_116; // @[Mem.scala 39:50:@1774.4]
  assign _T_1974 = io_mem_addr == 32'h75; // @[Mem.scala 39:41:@1781.4]
  assign _T_1975 = io_mem_wen & _T_1974; // @[Mem.scala 39:26:@1782.4]
  assign _GEN_15093 = _T_1975 ? io_mem_wdata : memory_117; // @[Mem.scala 39:50:@1783.4]
  assign _T_1983 = io_mem_addr == 32'h76; // @[Mem.scala 39:41:@1790.4]
  assign _T_1984 = io_mem_wen & _T_1983; // @[Mem.scala 39:26:@1791.4]
  assign _GEN_15222 = _T_1984 ? io_mem_wdata : memory_118; // @[Mem.scala 39:50:@1792.4]
  assign _T_1992 = io_mem_addr == 32'h77; // @[Mem.scala 39:41:@1799.4]
  assign _T_1993 = io_mem_wen & _T_1992; // @[Mem.scala 39:26:@1800.4]
  assign _GEN_15351 = _T_1993 ? io_mem_wdata : memory_119; // @[Mem.scala 39:50:@1801.4]
  assign _T_2001 = io_mem_addr == 32'h78; // @[Mem.scala 39:41:@1808.4]
  assign _T_2002 = io_mem_wen & _T_2001; // @[Mem.scala 39:26:@1809.4]
  assign _GEN_15480 = _T_2002 ? io_mem_wdata : memory_120; // @[Mem.scala 39:50:@1810.4]
  assign _T_2010 = io_mem_addr == 32'h79; // @[Mem.scala 39:41:@1817.4]
  assign _T_2011 = io_mem_wen & _T_2010; // @[Mem.scala 39:26:@1818.4]
  assign _GEN_15609 = _T_2011 ? io_mem_wdata : memory_121; // @[Mem.scala 39:50:@1819.4]
  assign _T_2019 = io_mem_addr == 32'h7a; // @[Mem.scala 39:41:@1826.4]
  assign _T_2020 = io_mem_wen & _T_2019; // @[Mem.scala 39:26:@1827.4]
  assign _GEN_15738 = _T_2020 ? io_mem_wdata : memory_122; // @[Mem.scala 39:50:@1828.4]
  assign _T_2028 = io_mem_addr == 32'h7b; // @[Mem.scala 39:41:@1835.4]
  assign _T_2029 = io_mem_wen & _T_2028; // @[Mem.scala 39:26:@1836.4]
  assign _GEN_15867 = _T_2029 ? io_mem_wdata : memory_123; // @[Mem.scala 39:50:@1837.4]
  assign _T_2037 = io_mem_addr == 32'h7c; // @[Mem.scala 39:41:@1844.4]
  assign _T_2038 = io_mem_wen & _T_2037; // @[Mem.scala 39:26:@1845.4]
  assign _GEN_15996 = _T_2038 ? io_mem_wdata : memory_124; // @[Mem.scala 39:50:@1846.4]
  assign _T_2046 = io_mem_addr == 32'h7d; // @[Mem.scala 39:41:@1853.4]
  assign _T_2047 = io_mem_wen & _T_2046; // @[Mem.scala 39:26:@1854.4]
  assign _GEN_16125 = _T_2047 ? io_mem_wdata : memory_125; // @[Mem.scala 39:50:@1855.4]
  assign _T_2055 = io_mem_addr == 32'h7e; // @[Mem.scala 39:41:@1862.4]
  assign _T_2056 = io_mem_wen & _T_2055; // @[Mem.scala 39:26:@1863.4]
  assign _GEN_16254 = _T_2056 ? io_mem_wdata : memory_126; // @[Mem.scala 39:50:@1864.4]
  assign _T_2064 = io_mem_addr == 32'h7f; // @[Mem.scala 39:41:@1871.4]
  assign _T_2065 = io_mem_wen & _T_2064; // @[Mem.scala 39:26:@1872.4]
  assign _GEN_16383 = _T_2065 ? io_mem_wdata : memory_127; // @[Mem.scala 39:50:@1873.4]
  assign io_mem_rdata = _T_2071; // @[Mem.scala 43:22:@736.4 Mem.scala 43:22:@745.4 Mem.scala 43:22:@754.4 Mem.scala 43:22:@763.4 Mem.scala 43:22:@772.4 Mem.scala 43:22:@781.4 Mem.scala 43:22:@790.4 Mem.scala 43:22:@799.4 Mem.scala 43:22:@808.4 Mem.scala 43:22:@817.4 Mem.scala 43:22:@826.4 Mem.scala 43:22:@835.4 Mem.scala 43:22:@844.4 Mem.scala 43:22:@853.4 Mem.scala 43:22:@862.4 Mem.scala 43:22:@871.4 Mem.scala 43:22:@880.4 Mem.scala 43:22:@889.4 Mem.scala 43:22:@898.4 Mem.scala 43:22:@907.4 Mem.scala 43:22:@916.4 Mem.scala 43:22:@925.4 Mem.scala 43:22:@934.4 Mem.scala 43:22:@943.4 Mem.scala 43:22:@952.4 Mem.scala 43:22:@961.4 Mem.scala 43:22:@970.4 Mem.scala 43:22:@979.4 Mem.scala 43:22:@988.4 Mem.scala 43:22:@997.4 Mem.scala 43:22:@1006.4 Mem.scala 43:22:@1015.4 Mem.scala 43:22:@1024.4 Mem.scala 43:22:@1033.4 Mem.scala 43:22:@1042.4 Mem.scala 43:22:@1051.4 Mem.scala 43:22:@1060.4 Mem.scala 43:22:@1069.4 Mem.scala 43:22:@1078.4 Mem.scala 43:22:@1087.4 Mem.scala 43:22:@1096.4 Mem.scala 43:22:@1105.4 Mem.scala 43:22:@1114.4 Mem.scala 43:22:@1123.4 Mem.scala 43:22:@1132.4 Mem.scala 43:22:@1141.4 Mem.scala 43:22:@1150.4 Mem.scala 43:22:@1159.4 Mem.scala 43:22:@1168.4 Mem.scala 43:22:@1177.4 Mem.scala 43:22:@1186.4 Mem.scala 43:22:@1195.4 Mem.scala 43:22:@1204.4 Mem.scala 43:22:@1213.4 Mem.scala 43:22:@1222.4 Mem.scala 43:22:@1231.4 Mem.scala 43:22:@1240.4 Mem.scala 43:22:@1249.4 Mem.scala 43:22:@1258.4 Mem.scala 43:22:@1267.4 Mem.scala 43:22:@1276.4 Mem.scala 43:22:@1285.4 Mem.scala 43:22:@1294.4 Mem.scala 43:22:@1303.4 Mem.scala 43:22:@1312.4 Mem.scala 43:22:@1321.4 Mem.scala 43:22:@1330.4 Mem.scala 43:22:@1339.4 Mem.scala 43:22:@1348.4 Mem.scala 43:22:@1357.4 Mem.scala 43:22:@1366.4 Mem.scala 43:22:@1375.4 Mem.scala 43:22:@1384.4 Mem.scala 43:22:@1393.4 Mem.scala 43:22:@1402.4 Mem.scala 43:22:@1411.4 Mem.scala 43:22:@1420.4 Mem.scala 43:22:@1429.4 Mem.scala 43:22:@1438.4 Mem.scala 43:22:@1447.4 Mem.scala 43:22:@1456.4 Mem.scala 43:22:@1465.4 Mem.scala 43:22:@1474.4 Mem.scala 43:22:@1483.4 Mem.scala 43:22:@1492.4 Mem.scala 43:22:@1501.4 Mem.scala 43:22:@1510.4 Mem.scala 43:22:@1519.4 Mem.scala 43:22:@1528.4 Mem.scala 43:22:@1537.4 Mem.scala 43:22:@1546.4 Mem.scala 43:22:@1555.4 Mem.scala 43:22:@1564.4 Mem.scala 43:22:@1573.4 Mem.scala 43:22:@1582.4 Mem.scala 43:22:@1591.4 Mem.scala 43:22:@1600.4 Mem.scala 43:22:@1609.4 Mem.scala 43:22:@1618.4 Mem.scala 43:22:@1627.4 Mem.scala 43:22:@1636.4 Mem.scala 43:22:@1645.4 Mem.scala 43:22:@1654.4 Mem.scala 43:22:@1663.4 Mem.scala 43:22:@1672.4 Mem.scala 43:22:@1681.4 Mem.scala 43:22:@1690.4 Mem.scala 43:22:@1699.4 Mem.scala 43:22:@1708.4 Mem.scala 43:22:@1717.4 Mem.scala 43:22:@1726.4 Mem.scala 43:22:@1735.4 Mem.scala 43:22:@1744.4 Mem.scala 43:22:@1753.4 Mem.scala 43:22:@1762.4 Mem.scala 43:22:@1771.4 Mem.scala 43:22:@1780.4 Mem.scala 43:22:@1789.4 Mem.scala 43:22:@1798.4 Mem.scala 43:22:@1807.4 Mem.scala 43:22:@1816.4 Mem.scala 43:22:@1825.4 Mem.scala 43:22:@1834.4 Mem.scala 43:22:@1843.4 Mem.scala 43:22:@1852.4 Mem.scala 43:22:@1861.4 Mem.scala 43:22:@1870.4 Mem.scala 43:22:@1879.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  memory_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  memory_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  memory_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  memory_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  memory_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  memory_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  memory_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  memory_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  memory_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  memory_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  memory_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  memory_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  memory_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  memory_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  memory_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  memory_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  memory_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  memory_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  memory_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  memory_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  memory_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  memory_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  memory_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  memory_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  memory_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  memory_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  memory_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  memory_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  memory_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  memory_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  memory_30 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  memory_31 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  memory_32 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  memory_33 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  memory_34 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  memory_35 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  memory_36 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  memory_37 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  memory_38 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  memory_39 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  memory_40 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  memory_41 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  memory_42 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  memory_43 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  memory_44 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  memory_45 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  memory_46 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  memory_47 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  memory_48 = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  memory_49 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  memory_50 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  memory_51 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  memory_52 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  memory_53 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  memory_54 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  memory_55 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  memory_56 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  memory_57 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  memory_58 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  memory_59 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  memory_60 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  memory_61 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  memory_62 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  memory_63 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  memory_64 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  memory_65 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  memory_66 = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  memory_67 = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  memory_68 = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  memory_69 = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  memory_70 = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  memory_71 = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  memory_72 = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  memory_73 = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  memory_74 = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  memory_75 = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  memory_76 = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  memory_77 = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  memory_78 = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  memory_79 = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  memory_80 = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  memory_81 = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  memory_82 = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  memory_83 = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  memory_84 = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  memory_85 = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  memory_86 = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  memory_87 = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  memory_88 = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  memory_89 = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  memory_90 = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  memory_91 = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  memory_92 = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  memory_93 = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  memory_94 = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  memory_95 = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  memory_96 = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  memory_97 = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  memory_98 = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  memory_99 = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  memory_100 = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  memory_101 = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  memory_102 = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  memory_103 = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  memory_104 = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  memory_105 = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  memory_106 = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  memory_107 = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  memory_108 = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  memory_109 = _RAND_109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  memory_110 = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  memory_111 = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  memory_112 = _RAND_112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  memory_113 = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  memory_114 = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  memory_115 = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  memory_116 = _RAND_116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  memory_117 = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  memory_118 = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  memory_119 = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  memory_120 = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  memory_121 = _RAND_121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  memory_122 = _RAND_122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  memory_123 = _RAND_123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  memory_124 = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  memory_125 = _RAND_125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  memory_126 = _RAND_126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  memory_127 = _RAND_127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_2071 = _RAND_128[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      memory_0 <= 32'h20010001;
    end else begin
      if (_T_922) begin
        memory_0 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_1 <= 32'h20210001;
    end else begin
      if (_T_931) begin
        memory_1 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_2 <= 32'h210820;
    end else begin
      if (_T_940) begin
        memory_2 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_3 <= 32'h8000002;
    end else begin
      if (_T_949) begin
        memory_3 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_4 <= 32'h8000003;
    end else begin
      if (_T_958) begin
        memory_4 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_5 <= 32'h8000003;
    end else begin
      if (_T_967) begin
        memory_5 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_6 <= 32'h8000003;
    end else begin
      if (_T_976) begin
        memory_6 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_7 <= 32'h8000003;
    end else begin
      if (_T_985) begin
        memory_7 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_8 <= 32'h0;
    end else begin
      if (_T_994) begin
        memory_8 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_9 <= 32'h0;
    end else begin
      if (_T_1003) begin
        memory_9 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_10 <= 32'h0;
    end else begin
      if (_T_1012) begin
        memory_10 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_11 <= 32'h0;
    end else begin
      if (_T_1021) begin
        memory_11 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_12 <= 32'h0;
    end else begin
      if (_T_1030) begin
        memory_12 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_13 <= 32'h0;
    end else begin
      if (_T_1039) begin
        memory_13 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_14 <= 32'h0;
    end else begin
      if (_T_1048) begin
        memory_14 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_15 <= 32'h0;
    end else begin
      if (_T_1057) begin
        memory_15 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_16 <= 32'h0;
    end else begin
      if (_T_1066) begin
        memory_16 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_17 <= 32'h0;
    end else begin
      if (_T_1075) begin
        memory_17 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_18 <= 32'h0;
    end else begin
      if (_T_1084) begin
        memory_18 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_19 <= 32'h0;
    end else begin
      if (_T_1093) begin
        memory_19 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_20 <= 32'h0;
    end else begin
      if (_T_1102) begin
        memory_20 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_21 <= 32'h0;
    end else begin
      if (_T_1111) begin
        memory_21 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_22 <= 32'h0;
    end else begin
      if (_T_1120) begin
        memory_22 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_23 <= 32'h0;
    end else begin
      if (_T_1129) begin
        memory_23 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_24 <= 32'h0;
    end else begin
      if (_T_1138) begin
        memory_24 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_25 <= 32'h0;
    end else begin
      if (_T_1147) begin
        memory_25 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_26 <= 32'h0;
    end else begin
      if (_T_1156) begin
        memory_26 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_27 <= 32'h0;
    end else begin
      if (_T_1165) begin
        memory_27 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_28 <= 32'h0;
    end else begin
      if (_T_1174) begin
        memory_28 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_29 <= 32'h0;
    end else begin
      if (_T_1183) begin
        memory_29 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_30 <= 32'h0;
    end else begin
      if (_T_1192) begin
        memory_30 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_31 <= 32'h0;
    end else begin
      if (_T_1201) begin
        memory_31 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_32 <= 32'h0;
    end else begin
      if (_T_1210) begin
        memory_32 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_33 <= 32'h0;
    end else begin
      if (_T_1219) begin
        memory_33 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_34 <= 32'h0;
    end else begin
      if (_T_1228) begin
        memory_34 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_35 <= 32'h0;
    end else begin
      if (_T_1237) begin
        memory_35 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_36 <= 32'h0;
    end else begin
      if (_T_1246) begin
        memory_36 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_37 <= 32'h0;
    end else begin
      if (_T_1255) begin
        memory_37 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_38 <= 32'h0;
    end else begin
      if (_T_1264) begin
        memory_38 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_39 <= 32'h0;
    end else begin
      if (_T_1273) begin
        memory_39 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_40 <= 32'h0;
    end else begin
      if (_T_1282) begin
        memory_40 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_41 <= 32'h0;
    end else begin
      if (_T_1291) begin
        memory_41 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_42 <= 32'h0;
    end else begin
      if (_T_1300) begin
        memory_42 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_43 <= 32'h0;
    end else begin
      if (_T_1309) begin
        memory_43 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_44 <= 32'h0;
    end else begin
      if (_T_1318) begin
        memory_44 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_45 <= 32'h0;
    end else begin
      if (_T_1327) begin
        memory_45 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_46 <= 32'h0;
    end else begin
      if (_T_1336) begin
        memory_46 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_47 <= 32'h0;
    end else begin
      if (_T_1345) begin
        memory_47 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_48 <= 32'h0;
    end else begin
      if (_T_1354) begin
        memory_48 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_49 <= 32'h0;
    end else begin
      if (_T_1363) begin
        memory_49 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_50 <= 32'h0;
    end else begin
      if (_T_1372) begin
        memory_50 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_51 <= 32'h0;
    end else begin
      if (_T_1381) begin
        memory_51 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_52 <= 32'h0;
    end else begin
      if (_T_1390) begin
        memory_52 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_53 <= 32'h0;
    end else begin
      if (_T_1399) begin
        memory_53 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_54 <= 32'h0;
    end else begin
      if (_T_1408) begin
        memory_54 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_55 <= 32'h0;
    end else begin
      if (_T_1417) begin
        memory_55 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_56 <= 32'h0;
    end else begin
      if (_T_1426) begin
        memory_56 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_57 <= 32'h0;
    end else begin
      if (_T_1435) begin
        memory_57 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_58 <= 32'h0;
    end else begin
      if (_T_1444) begin
        memory_58 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_59 <= 32'h0;
    end else begin
      if (_T_1453) begin
        memory_59 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_60 <= 32'h0;
    end else begin
      if (_T_1462) begin
        memory_60 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_61 <= 32'h0;
    end else begin
      if (_T_1471) begin
        memory_61 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_62 <= 32'h0;
    end else begin
      if (_T_1480) begin
        memory_62 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_63 <= 32'h0;
    end else begin
      if (_T_1489) begin
        memory_63 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_64 <= 32'h0;
    end else begin
      if (_T_1498) begin
        memory_64 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_65 <= 32'h0;
    end else begin
      if (_T_1507) begin
        memory_65 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_66 <= 32'h0;
    end else begin
      if (_T_1516) begin
        memory_66 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_67 <= 32'h0;
    end else begin
      if (_T_1525) begin
        memory_67 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_68 <= 32'h0;
    end else begin
      if (_T_1534) begin
        memory_68 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_69 <= 32'h0;
    end else begin
      if (_T_1543) begin
        memory_69 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_70 <= 32'h0;
    end else begin
      if (_T_1552) begin
        memory_70 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_71 <= 32'h0;
    end else begin
      if (_T_1561) begin
        memory_71 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_72 <= 32'h0;
    end else begin
      if (_T_1570) begin
        memory_72 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_73 <= 32'h0;
    end else begin
      if (_T_1579) begin
        memory_73 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_74 <= 32'h0;
    end else begin
      if (_T_1588) begin
        memory_74 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_75 <= 32'h0;
    end else begin
      if (_T_1597) begin
        memory_75 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_76 <= 32'h0;
    end else begin
      if (_T_1606) begin
        memory_76 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_77 <= 32'h0;
    end else begin
      if (_T_1615) begin
        memory_77 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_78 <= 32'h0;
    end else begin
      if (_T_1624) begin
        memory_78 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_79 <= 32'h0;
    end else begin
      if (_T_1633) begin
        memory_79 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_80 <= 32'h0;
    end else begin
      if (_T_1642) begin
        memory_80 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_81 <= 32'h0;
    end else begin
      if (_T_1651) begin
        memory_81 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_82 <= 32'h0;
    end else begin
      if (_T_1660) begin
        memory_82 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_83 <= 32'h0;
    end else begin
      if (_T_1669) begin
        memory_83 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_84 <= 32'h0;
    end else begin
      if (_T_1678) begin
        memory_84 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_85 <= 32'h0;
    end else begin
      if (_T_1687) begin
        memory_85 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_86 <= 32'h0;
    end else begin
      if (_T_1696) begin
        memory_86 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_87 <= 32'h0;
    end else begin
      if (_T_1705) begin
        memory_87 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_88 <= 32'h0;
    end else begin
      if (_T_1714) begin
        memory_88 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_89 <= 32'h0;
    end else begin
      if (_T_1723) begin
        memory_89 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_90 <= 32'h0;
    end else begin
      if (_T_1732) begin
        memory_90 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_91 <= 32'h0;
    end else begin
      if (_T_1741) begin
        memory_91 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_92 <= 32'h0;
    end else begin
      if (_T_1750) begin
        memory_92 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_93 <= 32'h0;
    end else begin
      if (_T_1759) begin
        memory_93 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_94 <= 32'h0;
    end else begin
      if (_T_1768) begin
        memory_94 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_95 <= 32'h0;
    end else begin
      if (_T_1777) begin
        memory_95 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_96 <= 32'h0;
    end else begin
      if (_T_1786) begin
        memory_96 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_97 <= 32'h0;
    end else begin
      if (_T_1795) begin
        memory_97 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_98 <= 32'h0;
    end else begin
      if (_T_1804) begin
        memory_98 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_99 <= 32'h0;
    end else begin
      if (_T_1813) begin
        memory_99 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_100 <= 32'h0;
    end else begin
      if (_T_1822) begin
        memory_100 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_101 <= 32'h0;
    end else begin
      if (_T_1831) begin
        memory_101 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_102 <= 32'h0;
    end else begin
      if (_T_1840) begin
        memory_102 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_103 <= 32'h0;
    end else begin
      if (_T_1849) begin
        memory_103 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_104 <= 32'h0;
    end else begin
      if (_T_1858) begin
        memory_104 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_105 <= 32'h0;
    end else begin
      if (_T_1867) begin
        memory_105 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_106 <= 32'h0;
    end else begin
      if (_T_1876) begin
        memory_106 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_107 <= 32'h0;
    end else begin
      if (_T_1885) begin
        memory_107 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_108 <= 32'h0;
    end else begin
      if (_T_1894) begin
        memory_108 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_109 <= 32'h0;
    end else begin
      if (_T_1903) begin
        memory_109 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_110 <= 32'h0;
    end else begin
      if (_T_1912) begin
        memory_110 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_111 <= 32'h0;
    end else begin
      if (_T_1921) begin
        memory_111 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_112 <= 32'h0;
    end else begin
      if (_T_1930) begin
        memory_112 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_113 <= 32'h0;
    end else begin
      if (_T_1939) begin
        memory_113 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_114 <= 32'h0;
    end else begin
      if (_T_1948) begin
        memory_114 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_115 <= 32'h0;
    end else begin
      if (_T_1957) begin
        memory_115 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_116 <= 32'h0;
    end else begin
      if (_T_1966) begin
        memory_116 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_117 <= 32'h0;
    end else begin
      if (_T_1975) begin
        memory_117 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_118 <= 32'h0;
    end else begin
      if (_T_1984) begin
        memory_118 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_119 <= 32'h0;
    end else begin
      if (_T_1993) begin
        memory_119 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_120 <= 32'h0;
    end else begin
      if (_T_2002) begin
        memory_120 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_121 <= 32'h0;
    end else begin
      if (_T_2011) begin
        memory_121 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_122 <= 32'h0;
    end else begin
      if (_T_2020) begin
        memory_122 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_123 <= 32'h0;
    end else begin
      if (_T_2029) begin
        memory_123 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_124 <= 32'h0;
    end else begin
      if (_T_2038) begin
        memory_124 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_125 <= 32'h0;
    end else begin
      if (_T_2047) begin
        memory_125 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_126 <= 32'h0;
    end else begin
      if (_T_2056) begin
        memory_126 <= io_mem_wdata;
      end
    end
    if (reset) begin
      memory_127 <= 32'h0;
    end else begin
      if (_T_2065) begin
        memory_127 <= io_mem_wdata;
      end
    end
    if (7'h7f == _T_926) begin
      _T_2071 <= memory_127;
    end else begin
      if (7'h7e == _T_926) begin
        _T_2071 <= memory_126;
      end else begin
        if (7'h7d == _T_926) begin
          _T_2071 <= memory_125;
        end else begin
          if (7'h7c == _T_926) begin
            _T_2071 <= memory_124;
          end else begin
            if (7'h7b == _T_926) begin
              _T_2071 <= memory_123;
            end else begin
              if (7'h7a == _T_926) begin
                _T_2071 <= memory_122;
              end else begin
                if (7'h79 == _T_926) begin
                  _T_2071 <= memory_121;
                end else begin
                  if (7'h78 == _T_926) begin
                    _T_2071 <= memory_120;
                  end else begin
                    if (7'h77 == _T_926) begin
                      _T_2071 <= memory_119;
                    end else begin
                      if (7'h76 == _T_926) begin
                        _T_2071 <= memory_118;
                      end else begin
                        if (7'h75 == _T_926) begin
                          _T_2071 <= memory_117;
                        end else begin
                          if (7'h74 == _T_926) begin
                            _T_2071 <= memory_116;
                          end else begin
                            if (7'h73 == _T_926) begin
                              _T_2071 <= memory_115;
                            end else begin
                              if (7'h72 == _T_926) begin
                                _T_2071 <= memory_114;
                              end else begin
                                if (7'h71 == _T_926) begin
                                  _T_2071 <= memory_113;
                                end else begin
                                  if (7'h70 == _T_926) begin
                                    _T_2071 <= memory_112;
                                  end else begin
                                    if (7'h6f == _T_926) begin
                                      _T_2071 <= memory_111;
                                    end else begin
                                      if (7'h6e == _T_926) begin
                                        _T_2071 <= memory_110;
                                      end else begin
                                        if (7'h6d == _T_926) begin
                                          _T_2071 <= memory_109;
                                        end else begin
                                          if (7'h6c == _T_926) begin
                                            _T_2071 <= memory_108;
                                          end else begin
                                            if (7'h6b == _T_926) begin
                                              _T_2071 <= memory_107;
                                            end else begin
                                              if (7'h6a == _T_926) begin
                                                _T_2071 <= memory_106;
                                              end else begin
                                                if (7'h69 == _T_926) begin
                                                  _T_2071 <= memory_105;
                                                end else begin
                                                  if (7'h68 == _T_926) begin
                                                    _T_2071 <= memory_104;
                                                  end else begin
                                                    if (7'h67 == _T_926) begin
                                                      _T_2071 <= memory_103;
                                                    end else begin
                                                      if (7'h66 == _T_926) begin
                                                        _T_2071 <= memory_102;
                                                      end else begin
                                                        if (7'h65 == _T_926) begin
                                                          _T_2071 <= memory_101;
                                                        end else begin
                                                          if (7'h64 == _T_926) begin
                                                            _T_2071 <= memory_100;
                                                          end else begin
                                                            if (7'h63 == _T_926) begin
                                                              _T_2071 <= memory_99;
                                                            end else begin
                                                              if (7'h62 == _T_926) begin
                                                                _T_2071 <= memory_98;
                                                              end else begin
                                                                if (7'h61 == _T_926) begin
                                                                  _T_2071 <= memory_97;
                                                                end else begin
                                                                  if (7'h60 == _T_926) begin
                                                                    _T_2071 <= memory_96;
                                                                  end else begin
                                                                    if (7'h5f == _T_926) begin
                                                                      _T_2071 <= memory_95;
                                                                    end else begin
                                                                      if (7'h5e == _T_926) begin
                                                                        _T_2071 <= memory_94;
                                                                      end else begin
                                                                        if (7'h5d == _T_926) begin
                                                                          _T_2071 <= memory_93;
                                                                        end else begin
                                                                          if (7'h5c == _T_926) begin
                                                                            _T_2071 <= memory_92;
                                                                          end else begin
                                                                            if (7'h5b == _T_926) begin
                                                                              _T_2071 <= memory_91;
                                                                            end else begin
                                                                              if (7'h5a == _T_926) begin
                                                                                _T_2071 <= memory_90;
                                                                              end else begin
                                                                                if (7'h59 == _T_926) begin
                                                                                  _T_2071 <= memory_89;
                                                                                end else begin
                                                                                  if (7'h58 == _T_926) begin
                                                                                    _T_2071 <= memory_88;
                                                                                  end else begin
                                                                                    if (7'h57 == _T_926) begin
                                                                                      _T_2071 <= memory_87;
                                                                                    end else begin
                                                                                      if (7'h56 == _T_926) begin
                                                                                        _T_2071 <= memory_86;
                                                                                      end else begin
                                                                                        if (7'h55 == _T_926) begin
                                                                                          _T_2071 <= memory_85;
                                                                                        end else begin
                                                                                          if (7'h54 == _T_926) begin
                                                                                            _T_2071 <= memory_84;
                                                                                          end else begin
                                                                                            if (7'h53 == _T_926) begin
                                                                                              _T_2071 <= memory_83;
                                                                                            end else begin
                                                                                              if (7'h52 == _T_926) begin
                                                                                                _T_2071 <= memory_82;
                                                                                              end else begin
                                                                                                if (7'h51 == _T_926) begin
                                                                                                  _T_2071 <= memory_81;
                                                                                                end else begin
                                                                                                  if (7'h50 == _T_926) begin
                                                                                                    _T_2071 <= memory_80;
                                                                                                  end else begin
                                                                                                    if (7'h4f == _T_926) begin
                                                                                                      _T_2071 <= memory_79;
                                                                                                    end else begin
                                                                                                      if (7'h4e == _T_926) begin
                                                                                                        _T_2071 <= memory_78;
                                                                                                      end else begin
                                                                                                        if (7'h4d == _T_926) begin
                                                                                                          _T_2071 <= memory_77;
                                                                                                        end else begin
                                                                                                          if (7'h4c == _T_926) begin
                                                                                                            _T_2071 <= memory_76;
                                                                                                          end else begin
                                                                                                            if (7'h4b == _T_926) begin
                                                                                                              _T_2071 <= memory_75;
                                                                                                            end else begin
                                                                                                              if (7'h4a == _T_926) begin
                                                                                                                _T_2071 <= memory_74;
                                                                                                              end else begin
                                                                                                                if (7'h49 == _T_926) begin
                                                                                                                  _T_2071 <= memory_73;
                                                                                                                end else begin
                                                                                                                  if (7'h48 == _T_926) begin
                                                                                                                    _T_2071 <= memory_72;
                                                                                                                  end else begin
                                                                                                                    if (7'h47 == _T_926) begin
                                                                                                                      _T_2071 <= memory_71;
                                                                                                                    end else begin
                                                                                                                      if (7'h46 == _T_926) begin
                                                                                                                        _T_2071 <= memory_70;
                                                                                                                      end else begin
                                                                                                                        if (7'h45 == _T_926) begin
                                                                                                                          _T_2071 <= memory_69;
                                                                                                                        end else begin
                                                                                                                          if (7'h44 == _T_926) begin
                                                                                                                            _T_2071 <= memory_68;
                                                                                                                          end else begin
                                                                                                                            if (7'h43 == _T_926) begin
                                                                                                                              _T_2071 <= memory_67;
                                                                                                                            end else begin
                                                                                                                              if (7'h42 == _T_926) begin
                                                                                                                                _T_2071 <= memory_66;
                                                                                                                              end else begin
                                                                                                                                if (7'h41 == _T_926) begin
                                                                                                                                  _T_2071 <= memory_65;
                                                                                                                                end else begin
                                                                                                                                  if (7'h40 == _T_926) begin
                                                                                                                                    _T_2071 <= memory_64;
                                                                                                                                  end else begin
                                                                                                                                    if (7'h3f == _T_926) begin
                                                                                                                                      _T_2071 <= memory_63;
                                                                                                                                    end else begin
                                                                                                                                      if (7'h3e == _T_926) begin
                                                                                                                                        _T_2071 <= memory_62;
                                                                                                                                      end else begin
                                                                                                                                        if (7'h3d == _T_926) begin
                                                                                                                                          _T_2071 <= memory_61;
                                                                                                                                        end else begin
                                                                                                                                          if (7'h3c == _T_926) begin
                                                                                                                                            _T_2071 <= memory_60;
                                                                                                                                          end else begin
                                                                                                                                            if (7'h3b == _T_926) begin
                                                                                                                                              _T_2071 <= memory_59;
                                                                                                                                            end else begin
                                                                                                                                              if (7'h3a == _T_926) begin
                                                                                                                                                _T_2071 <= memory_58;
                                                                                                                                              end else begin
                                                                                                                                                if (7'h39 == _T_926) begin
                                                                                                                                                  _T_2071 <= memory_57;
                                                                                                                                                end else begin
                                                                                                                                                  if (7'h38 == _T_926) begin
                                                                                                                                                    _T_2071 <= memory_56;
                                                                                                                                                  end else begin
                                                                                                                                                    if (7'h37 == _T_926) begin
                                                                                                                                                      _T_2071 <= memory_55;
                                                                                                                                                    end else begin
                                                                                                                                                      if (7'h36 == _T_926) begin
                                                                                                                                                        _T_2071 <= memory_54;
                                                                                                                                                      end else begin
                                                                                                                                                        if (7'h35 == _T_926) begin
                                                                                                                                                          _T_2071 <= memory_53;
                                                                                                                                                        end else begin
                                                                                                                                                          if (7'h34 == _T_926) begin
                                                                                                                                                            _T_2071 <= memory_52;
                                                                                                                                                          end else begin
                                                                                                                                                            if (7'h33 == _T_926) begin
                                                                                                                                                              _T_2071 <= memory_51;
                                                                                                                                                            end else begin
                                                                                                                                                              if (7'h32 == _T_926) begin
                                                                                                                                                                _T_2071 <= memory_50;
                                                                                                                                                              end else begin
                                                                                                                                                                if (7'h31 == _T_926) begin
                                                                                                                                                                  _T_2071 <= memory_49;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (7'h30 == _T_926) begin
                                                                                                                                                                    _T_2071 <= memory_48;
                                                                                                                                                                  end else begin
                                                                                                                                                                    if (7'h2f == _T_926) begin
                                                                                                                                                                      _T_2071 <= memory_47;
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (7'h2e == _T_926) begin
                                                                                                                                                                        _T_2071 <= memory_46;
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (7'h2d == _T_926) begin
                                                                                                                                                                          _T_2071 <= memory_45;
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (7'h2c == _T_926) begin
                                                                                                                                                                            _T_2071 <= memory_44;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (7'h2b == _T_926) begin
                                                                                                                                                                              _T_2071 <= memory_43;
                                                                                                                                                                            end else begin
                                                                                                                                                                              if (7'h2a == _T_926) begin
                                                                                                                                                                                _T_2071 <= memory_42;
                                                                                                                                                                              end else begin
                                                                                                                                                                                if (7'h29 == _T_926) begin
                                                                                                                                                                                  _T_2071 <= memory_41;
                                                                                                                                                                                end else begin
                                                                                                                                                                                  if (7'h28 == _T_926) begin
                                                                                                                                                                                    _T_2071 <= memory_40;
                                                                                                                                                                                  end else begin
                                                                                                                                                                                    if (7'h27 == _T_926) begin
                                                                                                                                                                                      _T_2071 <= memory_39;
                                                                                                                                                                                    end else begin
                                                                                                                                                                                      if (7'h26 == _T_926) begin
                                                                                                                                                                                        _T_2071 <= memory_38;
                                                                                                                                                                                      end else begin
                                                                                                                                                                                        if (7'h25 == _T_926) begin
                                                                                                                                                                                          _T_2071 <= memory_37;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                          if (7'h24 == _T_926) begin
                                                                                                                                                                                            _T_2071 <= memory_36;
                                                                                                                                                                                          end else begin
                                                                                                                                                                                            if (7'h23 == _T_926) begin
                                                                                                                                                                                              _T_2071 <= memory_35;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                              if (7'h22 == _T_926) begin
                                                                                                                                                                                                _T_2071 <= memory_34;
                                                                                                                                                                                              end else begin
                                                                                                                                                                                                if (7'h21 == _T_926) begin
                                                                                                                                                                                                  _T_2071 <= memory_33;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                  if (7'h20 == _T_926) begin
                                                                                                                                                                                                    _T_2071 <= memory_32;
                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                    if (7'h1f == _T_926) begin
                                                                                                                                                                                                      _T_2071 <= memory_31;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                      if (7'h1e == _T_926) begin
                                                                                                                                                                                                        _T_2071 <= memory_30;
                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                        if (7'h1d == _T_926) begin
                                                                                                                                                                                                          _T_2071 <= memory_29;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                          if (7'h1c == _T_926) begin
                                                                                                                                                                                                            _T_2071 <= memory_28;
                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                            if (7'h1b == _T_926) begin
                                                                                                                                                                                                              _T_2071 <= memory_27;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                              if (7'h1a == _T_926) begin
                                                                                                                                                                                                                _T_2071 <= memory_26;
                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                if (7'h19 == _T_926) begin
                                                                                                                                                                                                                  _T_2071 <= memory_25;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                  if (7'h18 == _T_926) begin
                                                                                                                                                                                                                    _T_2071 <= memory_24;
                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                    if (7'h17 == _T_926) begin
                                                                                                                                                                                                                      _T_2071 <= memory_23;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                      if (7'h16 == _T_926) begin
                                                                                                                                                                                                                        _T_2071 <= memory_22;
                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                        if (7'h15 == _T_926) begin
                                                                                                                                                                                                                          _T_2071 <= memory_21;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                          if (7'h14 == _T_926) begin
                                                                                                                                                                                                                            _T_2071 <= memory_20;
                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                            if (7'h13 == _T_926) begin
                                                                                                                                                                                                                              _T_2071 <= memory_19;
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                              if (7'h12 == _T_926) begin
                                                                                                                                                                                                                                _T_2071 <= memory_18;
                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                if (7'h11 == _T_926) begin
                                                                                                                                                                                                                                  _T_2071 <= memory_17;
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                  if (7'h10 == _T_926) begin
                                                                                                                                                                                                                                    _T_2071 <= memory_16;
                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                    if (7'hf == _T_926) begin
                                                                                                                                                                                                                                      _T_2071 <= memory_15;
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                      if (7'he == _T_926) begin
                                                                                                                                                                                                                                        _T_2071 <= memory_14;
                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                        if (7'hd == _T_926) begin
                                                                                                                                                                                                                                          _T_2071 <= memory_13;
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                          if (7'hc == _T_926) begin
                                                                                                                                                                                                                                            _T_2071 <= memory_12;
                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                            if (7'hb == _T_926) begin
                                                                                                                                                                                                                                              _T_2071 <= memory_11;
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                              if (7'ha == _T_926) begin
                                                                                                                                                                                                                                                _T_2071 <= memory_10;
                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                if (7'h9 == _T_926) begin
                                                                                                                                                                                                                                                  _T_2071 <= memory_9;
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                  if (7'h8 == _T_926) begin
                                                                                                                                                                                                                                                    _T_2071 <= memory_8;
                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                    if (7'h7 == _T_926) begin
                                                                                                                                                                                                                                                      _T_2071 <= memory_7;
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                      if (7'h6 == _T_926) begin
                                                                                                                                                                                                                                                        _T_2071 <= memory_6;
                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                        if (7'h5 == _T_926) begin
                                                                                                                                                                                                                                                          _T_2071 <= memory_5;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                          if (7'h4 == _T_926) begin
                                                                                                                                                                                                                                                            _T_2071 <= memory_4;
                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                            if (7'h3 == _T_926) begin
                                                                                                                                                                                                                                                              _T_2071 <= memory_3;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                              if (7'h2 == _T_926) begin
                                                                                                                                                                                                                                                                _T_2071 <= memory_2;
                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                if (7'h1 == _T_926) begin
                                                                                                                                                                                                                                                                  _T_2071 <= memory_1;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                  _T_2071 <= memory_0;
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                              end
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                          end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                      end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                  end
                                                                                                                                                                                                                end
                                                                                                                                                                                                              end
                                                                                                                                                                                                            end
                                                                                                                                                                                                          end
                                                                                                                                                                                                        end
                                                                                                                                                                                                      end
                                                                                                                                                                                                    end
                                                                                                                                                                                                  end
                                                                                                                                                                                                end
                                                                                                                                                                                              end
                                                                                                                                                                                            end
                                                                                                                                                                                          end
                                                                                                                                                                                        end
                                                                                                                                                                                      end
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end
                                                                                                                                                      end
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end
                                                                                                                                        end
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module CPU( // @[:@1881.2]
  input         clock, // @[:@1882.4]
  input         reset, // @[:@1883.4]
  output [31:0] io_debug_ir, // @[:@1884.4]
  output [31:0] io_debug_mdr, // @[:@1884.4]
  output [31:0] io_debug_aluout, // @[:@1884.4]
  output [31:0] io_debug_pc, // @[:@1884.4]
  input  [4:0]  io_debug_ra_c, // @[:@1884.4]
  output [31:0] io_debug_rd_c, // @[:@1884.4]
  output [3:0]  io_ctrl_dbg_cur_state, // @[:@1884.4]
  output        io_ctrl_dbg_isRType, // @[:@1884.4]
  output        io_ctrl_dbg_isIType, // @[:@1884.4]
  output        io_ctrl_dbg_isJType, // @[:@1884.4]
  output        io_ctrl_dbg_isLW, // @[:@1884.4]
  output        io_ctrl_dbg_isSW, // @[:@1884.4]
  output        io_ctrl_dbg_isBEQ, // @[:@1884.4]
  output        io_ctrl_dbg_isBNE // @[:@1884.4]
);
  wire  datapath_clock; // @[CPU.scala 30:26:@1886.4]
  wire  datapath_reset; // @[CPU.scala 30:26:@1886.4]
  wire [31:0] datapath_io_ctrl_Inst; // @[CPU.scala 30:26:@1886.4]
  wire  datapath_io_ctrl_IRWrite; // @[CPU.scala 30:26:@1886.4]
  wire  datapath_io_ctrl_RegDst; // @[CPU.scala 30:26:@1886.4]
  wire  datapath_io_ctrl_RegWrite; // @[CPU.scala 30:26:@1886.4]
  wire  datapath_io_ctrl_ALUSrcA; // @[CPU.scala 30:26:@1886.4]
  wire [2:0] datapath_io_ctrl_ALUSrcB; // @[CPU.scala 30:26:@1886.4]
  wire [3:0] datapath_io_ctrl_ALUOp; // @[CPU.scala 30:26:@1886.4]
  wire [1:0] datapath_io_ctrl_PCSource; // @[CPU.scala 30:26:@1886.4]
  wire  datapath_io_ctrl_PCWriteBEQ; // @[CPU.scala 30:26:@1886.4]
  wire  datapath_io_ctrl_PCWriteBNE; // @[CPU.scala 30:26:@1886.4]
  wire  datapath_io_ctrl_PCWrite; // @[CPU.scala 30:26:@1886.4]
  wire  datapath_io_ctrl_IorD; // @[CPU.scala 30:26:@1886.4]
  wire  datapath_io_ctrl_MemWrite; // @[CPU.scala 30:26:@1886.4]
  wire  datapath_io_ctrl_MemtoReg; // @[CPU.scala 30:26:@1886.4]
  wire [31:0] datapath_io_mem_mem_rdata; // @[CPU.scala 30:26:@1886.4]
  wire [31:0] datapath_io_mem_mem_addr; // @[CPU.scala 30:26:@1886.4]
  wire [31:0] datapath_io_mem_mem_wdata; // @[CPU.scala 30:26:@1886.4]
  wire  datapath_io_mem_mem_wen; // @[CPU.scala 30:26:@1886.4]
  wire [31:0] datapath_io_debug_ir; // @[CPU.scala 30:26:@1886.4]
  wire [31:0] datapath_io_debug_mdr; // @[CPU.scala 30:26:@1886.4]
  wire [31:0] datapath_io_debug_aluout; // @[CPU.scala 30:26:@1886.4]
  wire [31:0] datapath_io_debug_pc; // @[CPU.scala 30:26:@1886.4]
  wire [4:0] datapath_io_debug_ra_c; // @[CPU.scala 30:26:@1886.4]
  wire [31:0] datapath_io_debug_rd_c; // @[CPU.scala 30:26:@1886.4]
  wire  ctrl_clock; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_reset; // @[CPU.scala 33:22:@1895.4]
  wire [31:0] ctrl_io_Inst; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_io_IRWrite; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_io_RegDst; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_io_RegWrite; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_io_ALUSrcA; // @[CPU.scala 33:22:@1895.4]
  wire [2:0] ctrl_io_ALUSrcB; // @[CPU.scala 33:22:@1895.4]
  wire [3:0] ctrl_io_ALUOp; // @[CPU.scala 33:22:@1895.4]
  wire [1:0] ctrl_io_PCSource; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_io_PCWriteBEQ; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_io_PCWriteBNE; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_io_PCWrite; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_io_IorD; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_io_MemWrite; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_io_MemtoReg; // @[CPU.scala 33:22:@1895.4]
  wire [3:0] ctrl_io_ctrl_dbg_cur_state; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_io_ctrl_dbg_isRType; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_io_ctrl_dbg_isIType; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_io_ctrl_dbg_isJType; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_io_ctrl_dbg_isLW; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_io_ctrl_dbg_isSW; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_io_ctrl_dbg_isBEQ; // @[CPU.scala 33:22:@1895.4]
  wire  ctrl_io_ctrl_dbg_isBNE; // @[CPU.scala 33:22:@1895.4]
  wire  mem_clock; // @[CPU.scala 37:21:@1929.4]
  wire  mem_reset; // @[CPU.scala 37:21:@1929.4]
  wire [31:0] mem_io_mem_rdata; // @[CPU.scala 37:21:@1929.4]
  wire [31:0] mem_io_mem_addr; // @[CPU.scala 37:21:@1929.4]
  wire [31:0] mem_io_mem_wdata; // @[CPU.scala 37:21:@1929.4]
  wire  mem_io_mem_wen; // @[CPU.scala 37:21:@1929.4]
  Datapath datapath ( // @[CPU.scala 30:26:@1886.4]
    .clock(datapath_clock),
    .reset(datapath_reset),
    .io_ctrl_Inst(datapath_io_ctrl_Inst),
    .io_ctrl_IRWrite(datapath_io_ctrl_IRWrite),
    .io_ctrl_RegDst(datapath_io_ctrl_RegDst),
    .io_ctrl_RegWrite(datapath_io_ctrl_RegWrite),
    .io_ctrl_ALUSrcA(datapath_io_ctrl_ALUSrcA),
    .io_ctrl_ALUSrcB(datapath_io_ctrl_ALUSrcB),
    .io_ctrl_ALUOp(datapath_io_ctrl_ALUOp),
    .io_ctrl_PCSource(datapath_io_ctrl_PCSource),
    .io_ctrl_PCWriteBEQ(datapath_io_ctrl_PCWriteBEQ),
    .io_ctrl_PCWriteBNE(datapath_io_ctrl_PCWriteBNE),
    .io_ctrl_PCWrite(datapath_io_ctrl_PCWrite),
    .io_ctrl_IorD(datapath_io_ctrl_IorD),
    .io_ctrl_MemWrite(datapath_io_ctrl_MemWrite),
    .io_ctrl_MemtoReg(datapath_io_ctrl_MemtoReg),
    .io_mem_mem_rdata(datapath_io_mem_mem_rdata),
    .io_mem_mem_addr(datapath_io_mem_mem_addr),
    .io_mem_mem_wdata(datapath_io_mem_mem_wdata),
    .io_mem_mem_wen(datapath_io_mem_mem_wen),
    .io_debug_ir(datapath_io_debug_ir),
    .io_debug_mdr(datapath_io_debug_mdr),
    .io_debug_aluout(datapath_io_debug_aluout),
    .io_debug_pc(datapath_io_debug_pc),
    .io_debug_ra_c(datapath_io_debug_ra_c),
    .io_debug_rd_c(datapath_io_debug_rd_c)
  );
  Control ctrl ( // @[CPU.scala 33:22:@1895.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_Inst(ctrl_io_Inst),
    .io_IRWrite(ctrl_io_IRWrite),
    .io_RegDst(ctrl_io_RegDst),
    .io_RegWrite(ctrl_io_RegWrite),
    .io_ALUSrcA(ctrl_io_ALUSrcA),
    .io_ALUSrcB(ctrl_io_ALUSrcB),
    .io_ALUOp(ctrl_io_ALUOp),
    .io_PCSource(ctrl_io_PCSource),
    .io_PCWriteBEQ(ctrl_io_PCWriteBEQ),
    .io_PCWriteBNE(ctrl_io_PCWriteBNE),
    .io_PCWrite(ctrl_io_PCWrite),
    .io_IorD(ctrl_io_IorD),
    .io_MemWrite(ctrl_io_MemWrite),
    .io_MemtoReg(ctrl_io_MemtoReg),
    .io_ctrl_dbg_cur_state(ctrl_io_ctrl_dbg_cur_state),
    .io_ctrl_dbg_isRType(ctrl_io_ctrl_dbg_isRType),
    .io_ctrl_dbg_isIType(ctrl_io_ctrl_dbg_isIType),
    .io_ctrl_dbg_isJType(ctrl_io_ctrl_dbg_isJType),
    .io_ctrl_dbg_isLW(ctrl_io_ctrl_dbg_isLW),
    .io_ctrl_dbg_isSW(ctrl_io_ctrl_dbg_isSW),
    .io_ctrl_dbg_isBEQ(ctrl_io_ctrl_dbg_isBEQ),
    .io_ctrl_dbg_isBNE(ctrl_io_ctrl_dbg_isBNE)
  );
  Mem mem ( // @[CPU.scala 37:21:@1929.4]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_mem_rdata(mem_io_mem_rdata),
    .io_mem_addr(mem_io_mem_addr),
    .io_mem_wdata(mem_io_mem_wdata),
    .io_mem_wen(mem_io_mem_wen)
  );
  assign io_debug_ir = datapath_io_debug_ir; // @[CPU.scala 31:14:@1894.4]
  assign io_debug_mdr = datapath_io_debug_mdr; // @[CPU.scala 31:14:@1893.4]
  assign io_debug_aluout = datapath_io_debug_aluout; // @[CPU.scala 31:14:@1892.4]
  assign io_debug_pc = datapath_io_debug_pc; // @[CPU.scala 31:14:@1891.4]
  assign io_debug_rd_c = datapath_io_debug_rd_c; // @[CPU.scala 31:14:@1889.4]
  assign io_ctrl_dbg_cur_state = ctrl_io_ctrl_dbg_cur_state; // @[CPU.scala 35:17:@1928.4]
  assign io_ctrl_dbg_isRType = ctrl_io_ctrl_dbg_isRType; // @[CPU.scala 35:17:@1927.4]
  assign io_ctrl_dbg_isIType = ctrl_io_ctrl_dbg_isIType; // @[CPU.scala 35:17:@1926.4]
  assign io_ctrl_dbg_isJType = ctrl_io_ctrl_dbg_isJType; // @[CPU.scala 35:17:@1925.4]
  assign io_ctrl_dbg_isLW = ctrl_io_ctrl_dbg_isLW; // @[CPU.scala 35:17:@1924.4]
  assign io_ctrl_dbg_isSW = ctrl_io_ctrl_dbg_isSW; // @[CPU.scala 35:17:@1923.4]
  assign io_ctrl_dbg_isBEQ = ctrl_io_ctrl_dbg_isBEQ; // @[CPU.scala 35:17:@1922.4]
  assign io_ctrl_dbg_isBNE = ctrl_io_ctrl_dbg_isBNE; // @[CPU.scala 35:17:@1921.4]
  assign datapath_clock = clock; // @[:@1887.4]
  assign datapath_reset = reset; // @[:@1888.4]
  assign datapath_io_ctrl_IRWrite = ctrl_io_IRWrite; // @[CPU.scala 34:13:@1919.4]
  assign datapath_io_ctrl_RegDst = ctrl_io_RegDst; // @[CPU.scala 34:13:@1918.4]
  assign datapath_io_ctrl_RegWrite = ctrl_io_RegWrite; // @[CPU.scala 34:13:@1917.4]
  assign datapath_io_ctrl_ALUSrcA = ctrl_io_ALUSrcA; // @[CPU.scala 34:13:@1916.4]
  assign datapath_io_ctrl_ALUSrcB = ctrl_io_ALUSrcB; // @[CPU.scala 34:13:@1915.4]
  assign datapath_io_ctrl_ALUOp = ctrl_io_ALUOp; // @[CPU.scala 34:13:@1914.4]
  assign datapath_io_ctrl_PCSource = ctrl_io_PCSource; // @[CPU.scala 34:13:@1913.4]
  assign datapath_io_ctrl_PCWriteBEQ = ctrl_io_PCWriteBEQ; // @[CPU.scala 34:13:@1912.4]
  assign datapath_io_ctrl_PCWriteBNE = ctrl_io_PCWriteBNE; // @[CPU.scala 34:13:@1911.4]
  assign datapath_io_ctrl_PCWrite = ctrl_io_PCWrite; // @[CPU.scala 34:13:@1910.4]
  assign datapath_io_ctrl_IorD = ctrl_io_IorD; // @[CPU.scala 34:13:@1909.4]
  assign datapath_io_ctrl_MemWrite = ctrl_io_MemWrite; // @[CPU.scala 34:13:@1907.4]
  assign datapath_io_ctrl_MemtoReg = ctrl_io_MemtoReg; // @[CPU.scala 34:13:@1906.4]
  assign datapath_io_mem_mem_rdata = mem_io_mem_rdata; // @[CPU.scala 38:12:@1935.4]
  assign datapath_io_debug_ra_c = io_debug_ra_c; // @[CPU.scala 31:14:@1890.4]
  assign ctrl_clock = clock; // @[:@1896.4]
  assign ctrl_reset = reset; // @[:@1897.4]
  assign ctrl_io_Inst = datapath_io_ctrl_Inst; // @[CPU.scala 34:13:@1920.4]
  assign mem_clock = clock; // @[:@1930.4]
  assign mem_reset = reset; // @[:@1931.4]
  assign mem_io_mem_addr = datapath_io_mem_mem_addr; // @[CPU.scala 38:12:@1934.4]
  assign mem_io_mem_wdata = datapath_io_mem_mem_wdata; // @[CPU.scala 38:12:@1933.4]
  assign mem_io_mem_wen = datapath_io_mem_mem_wen; // @[CPU.scala 38:12:@1932.4]
endmodule
