module ALU( // @[:@3.2]
  input  [31:0] io_A, // @[:@6.4]
  input  [31:0] io_B, // @[:@6.4]
  input  [3:0]  io_opcode, // @[:@6.4]
  output [31:0] io_out, // @[:@6.4]
  output        io_flagZero // @[:@6.4]
);
  wire [32:0] _T_29; // @[ALU.scala 34:32:@8.4]
  wire [31:0] _T_30; // @[ALU.scala 34:32:@9.4]
  wire [32:0] _T_31; // @[ALU.scala 35:32:@10.4]
  wire [32:0] _T_32; // @[ALU.scala 35:32:@11.4]
  wire [31:0] _T_33; // @[ALU.scala 35:32:@12.4]
  wire [4:0] _T_34; // @[ALU.scala 38:39:@13.4]
  wire [62:0] _GEN_0; // @[ALU.scala 38:32:@14.4]
  wire [62:0] _T_35; // @[ALU.scala 38:32:@14.4]
  wire [31:0] _T_36; // @[ALU.scala 39:32:@15.4]
  wire [31:0] _T_37; // @[ALU.scala 39:46:@16.4]
  wire  _T_38; // @[ALU.scala 39:39:@17.4]
  wire  _T_39; // @[ALU.scala 40:32:@18.4]
  wire [31:0] _T_40; // @[ALU.scala 41:32:@19.4]
  wire [31:0] _T_41; // @[ALU.scala 42:32:@20.4]
  wire [31:0] _T_42; // @[ALU.scala 43:32:@21.4]
  wire [31:0] _T_44; // @[ALU.scala 44:26:@23.4]
  wire  _T_45; // @[Mux.scala 46:19:@24.4]
  wire [31:0] _T_46; // @[Mux.scala 46:16:@25.4]
  wire  _T_47; // @[Mux.scala 46:19:@26.4]
  wire [31:0] _T_48; // @[Mux.scala 46:16:@27.4]
  wire  _T_49; // @[Mux.scala 46:19:@28.4]
  wire [31:0] _T_50; // @[Mux.scala 46:16:@29.4]
  wire  _T_51; // @[Mux.scala 46:19:@30.4]
  wire [31:0] _T_52; // @[Mux.scala 46:16:@31.4]
  wire  _T_53; // @[Mux.scala 46:19:@32.4]
  wire [31:0] _T_54; // @[Mux.scala 46:16:@33.4]
  wire  _T_55; // @[Mux.scala 46:19:@34.4]
  wire [31:0] _T_56; // @[Mux.scala 46:16:@35.4]
  wire  _T_57; // @[Mux.scala 46:19:@36.4]
  wire [31:0] _T_58; // @[Mux.scala 46:16:@37.4]
  wire  _T_59; // @[Mux.scala 46:19:@38.4]
  wire [62:0] _T_60; // @[Mux.scala 46:16:@39.4]
  wire  _T_61; // @[Mux.scala 46:19:@40.4]
  wire [62:0] _T_62; // @[Mux.scala 46:16:@41.4]
  wire  _T_63; // @[Mux.scala 46:19:@42.4]
  wire [62:0] _T_64; // @[Mux.scala 46:16:@43.4]
  assign _T_29 = io_A + io_B; // @[ALU.scala 34:32:@8.4]
  assign _T_30 = io_A + io_B; // @[ALU.scala 34:32:@9.4]
  assign _T_31 = io_A - io_B; // @[ALU.scala 35:32:@10.4]
  assign _T_32 = $unsigned(_T_31); // @[ALU.scala 35:32:@11.4]
  assign _T_33 = _T_32[31:0]; // @[ALU.scala 35:32:@12.4]
  assign _T_34 = io_B[4:0]; // @[ALU.scala 38:39:@13.4]
  assign _GEN_0 = {{31'd0}, io_A}; // @[ALU.scala 38:32:@14.4]
  assign _T_35 = _GEN_0 << _T_34; // @[ALU.scala 38:32:@14.4]
  assign _T_36 = $signed(io_A); // @[ALU.scala 39:32:@15.4]
  assign _T_37 = $signed(io_B); // @[ALU.scala 39:46:@16.4]
  assign _T_38 = $signed(_T_36) < $signed(_T_37); // @[ALU.scala 39:39:@17.4]
  assign _T_39 = io_A < io_B; // @[ALU.scala 40:32:@18.4]
  assign _T_40 = io_A & io_B; // @[ALU.scala 41:32:@19.4]
  assign _T_41 = io_A | io_B; // @[ALU.scala 42:32:@20.4]
  assign _T_42 = io_A ^ io_B; // @[ALU.scala 43:32:@21.4]
  assign _T_44 = ~ _T_41; // @[ALU.scala 44:26:@23.4]
  assign _T_45 = 4'ha == io_opcode; // @[Mux.scala 46:19:@24.4]
  assign _T_46 = _T_45 ? io_A : io_B; // @[Mux.scala 46:16:@25.4]
  assign _T_47 = 4'hc == io_opcode; // @[Mux.scala 46:19:@26.4]
  assign _T_48 = _T_47 ? _T_44 : _T_46; // @[Mux.scala 46:16:@27.4]
  assign _T_49 = 4'h4 == io_opcode; // @[Mux.scala 46:19:@28.4]
  assign _T_50 = _T_49 ? _T_42 : _T_48; // @[Mux.scala 46:16:@29.4]
  assign _T_51 = 4'h3 == io_opcode; // @[Mux.scala 46:19:@30.4]
  assign _T_52 = _T_51 ? _T_41 : _T_50; // @[Mux.scala 46:16:@31.4]
  assign _T_53 = 4'h2 == io_opcode; // @[Mux.scala 46:19:@32.4]
  assign _T_54 = _T_53 ? _T_40 : _T_52; // @[Mux.scala 46:16:@33.4]
  assign _T_55 = 4'h7 == io_opcode; // @[Mux.scala 46:19:@34.4]
  assign _T_56 = _T_55 ? {{31'd0}, _T_39} : _T_54; // @[Mux.scala 46:16:@35.4]
  assign _T_57 = 4'h5 == io_opcode; // @[Mux.scala 46:19:@36.4]
  assign _T_58 = _T_57 ? {{31'd0}, _T_38} : _T_56; // @[Mux.scala 46:16:@37.4]
  assign _T_59 = 4'h6 == io_opcode; // @[Mux.scala 46:19:@38.4]
  assign _T_60 = _T_59 ? _T_35 : {{31'd0}, _T_58}; // @[Mux.scala 46:16:@39.4]
  assign _T_61 = 4'h1 == io_opcode; // @[Mux.scala 46:19:@40.4]
  assign _T_62 = _T_61 ? {{31'd0}, _T_33} : _T_60; // @[Mux.scala 46:16:@41.4]
  assign _T_63 = 4'h0 == io_opcode; // @[Mux.scala 46:19:@42.4]
  assign _T_64 = _T_63 ? {{31'd0}, _T_30} : _T_62; // @[Mux.scala 46:16:@43.4]
  assign io_out = _T_64[31:0]; // @[ALU.scala 33:12:@44.4]
  assign io_flagZero = io_out == 32'h0; // @[ALU.scala 47:17:@46.4]
endmodule
module RegFile( // @[:@48.2]
  input         clock, // @[:@49.4]
  input         reset, // @[:@50.4]
  input  [4:0]  io_ra_a, // @[:@51.4]
  input  [4:0]  io_ra_b, // @[:@51.4]
  input  [4:0]  io_wa, // @[:@51.4]
  input  [31:0] io_wd, // @[:@51.4]
  output [31:0] io_rd_a, // @[:@51.4]
  output [31:0] io_rd_b, // @[:@51.4]
  input         io_RegWrite, // @[:@51.4]
  input  [4:0]  io_ra_c, // @[:@51.4]
  output [31:0] io_rd_c // @[:@51.4]
);
  reg [31:0] regs_0; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_0;
  reg [31:0] regs_1; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_1;
  reg [31:0] regs_2; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_2;
  reg [31:0] regs_3; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_3;
  reg [31:0] regs_4; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_4;
  reg [31:0] regs_5; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_5;
  reg [31:0] regs_6; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_6;
  reg [31:0] regs_7; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_7;
  reg [31:0] regs_8; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_8;
  reg [31:0] regs_9; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_9;
  reg [31:0] regs_10; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_10;
  reg [31:0] regs_11; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_11;
  reg [31:0] regs_12; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_12;
  reg [31:0] regs_13; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_13;
  reg [31:0] regs_14; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_14;
  reg [31:0] regs_15; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_15;
  reg [31:0] regs_16; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_16;
  reg [31:0] regs_17; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_17;
  reg [31:0] regs_18; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_18;
  reg [31:0] regs_19; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_19;
  reg [31:0] regs_20; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_20;
  reg [31:0] regs_21; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_21;
  reg [31:0] regs_22; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_22;
  reg [31:0] regs_23; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_23;
  reg [31:0] regs_24; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_24;
  reg [31:0] regs_25; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_25;
  reg [31:0] regs_26; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_26;
  reg [31:0] regs_27; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_27;
  reg [31:0] regs_28; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_28;
  reg [31:0] regs_29; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_29;
  reg [31:0] regs_30; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_30;
  reg [31:0] regs_31; // @[RegFile.scala 21:23:@86.4]
  reg [31:0] _RAND_31;
  wire  _T_262; // @[RegFile.scala 23:21:@87.4]
  wire  _T_263; // @[RegFile.scala 23:34:@88.4]
  wire [31:0] _GEN_0; // @[RegFile.scala 23:50:@89.4]
  wire  _T_265; // @[RegFile.scala 23:21:@92.4]
  wire  _T_266; // @[RegFile.scala 23:34:@93.4]
  wire [31:0] _GEN_1; // @[RegFile.scala 23:50:@94.4]
  wire  _T_268; // @[RegFile.scala 23:21:@97.4]
  wire  _T_269; // @[RegFile.scala 23:34:@98.4]
  wire [31:0] _GEN_2; // @[RegFile.scala 23:50:@99.4]
  wire  _T_271; // @[RegFile.scala 23:21:@102.4]
  wire  _T_272; // @[RegFile.scala 23:34:@103.4]
  wire [31:0] _GEN_3; // @[RegFile.scala 23:50:@104.4]
  wire  _T_274; // @[RegFile.scala 23:21:@107.4]
  wire  _T_275; // @[RegFile.scala 23:34:@108.4]
  wire [31:0] _GEN_4; // @[RegFile.scala 23:50:@109.4]
  wire  _T_277; // @[RegFile.scala 23:21:@112.4]
  wire  _T_278; // @[RegFile.scala 23:34:@113.4]
  wire [31:0] _GEN_5; // @[RegFile.scala 23:50:@114.4]
  wire  _T_280; // @[RegFile.scala 23:21:@117.4]
  wire  _T_281; // @[RegFile.scala 23:34:@118.4]
  wire [31:0] _GEN_6; // @[RegFile.scala 23:50:@119.4]
  wire  _T_283; // @[RegFile.scala 23:21:@122.4]
  wire  _T_284; // @[RegFile.scala 23:34:@123.4]
  wire [31:0] _GEN_7; // @[RegFile.scala 23:50:@124.4]
  wire  _T_286; // @[RegFile.scala 23:21:@127.4]
  wire  _T_287; // @[RegFile.scala 23:34:@128.4]
  wire [31:0] _GEN_8; // @[RegFile.scala 23:50:@129.4]
  wire  _T_289; // @[RegFile.scala 23:21:@132.4]
  wire  _T_290; // @[RegFile.scala 23:34:@133.4]
  wire [31:0] _GEN_9; // @[RegFile.scala 23:50:@134.4]
  wire  _T_292; // @[RegFile.scala 23:21:@137.4]
  wire  _T_293; // @[RegFile.scala 23:34:@138.4]
  wire [31:0] _GEN_10; // @[RegFile.scala 23:50:@139.4]
  wire  _T_295; // @[RegFile.scala 23:21:@142.4]
  wire  _T_296; // @[RegFile.scala 23:34:@143.4]
  wire [31:0] _GEN_11; // @[RegFile.scala 23:50:@144.4]
  wire  _T_298; // @[RegFile.scala 23:21:@147.4]
  wire  _T_299; // @[RegFile.scala 23:34:@148.4]
  wire [31:0] _GEN_12; // @[RegFile.scala 23:50:@149.4]
  wire  _T_301; // @[RegFile.scala 23:21:@152.4]
  wire  _T_302; // @[RegFile.scala 23:34:@153.4]
  wire [31:0] _GEN_13; // @[RegFile.scala 23:50:@154.4]
  wire  _T_304; // @[RegFile.scala 23:21:@157.4]
  wire  _T_305; // @[RegFile.scala 23:34:@158.4]
  wire [31:0] _GEN_14; // @[RegFile.scala 23:50:@159.4]
  wire  _T_307; // @[RegFile.scala 23:21:@162.4]
  wire  _T_308; // @[RegFile.scala 23:34:@163.4]
  wire [31:0] _GEN_15; // @[RegFile.scala 23:50:@164.4]
  wire  _T_310; // @[RegFile.scala 23:21:@167.4]
  wire  _T_311; // @[RegFile.scala 23:34:@168.4]
  wire [31:0] _GEN_16; // @[RegFile.scala 23:50:@169.4]
  wire  _T_313; // @[RegFile.scala 23:21:@172.4]
  wire  _T_314; // @[RegFile.scala 23:34:@173.4]
  wire [31:0] _GEN_17; // @[RegFile.scala 23:50:@174.4]
  wire  _T_316; // @[RegFile.scala 23:21:@177.4]
  wire  _T_317; // @[RegFile.scala 23:34:@178.4]
  wire [31:0] _GEN_18; // @[RegFile.scala 23:50:@179.4]
  wire  _T_319; // @[RegFile.scala 23:21:@182.4]
  wire  _T_320; // @[RegFile.scala 23:34:@183.4]
  wire [31:0] _GEN_19; // @[RegFile.scala 23:50:@184.4]
  wire  _T_322; // @[RegFile.scala 23:21:@187.4]
  wire  _T_323; // @[RegFile.scala 23:34:@188.4]
  wire [31:0] _GEN_20; // @[RegFile.scala 23:50:@189.4]
  wire  _T_325; // @[RegFile.scala 23:21:@192.4]
  wire  _T_326; // @[RegFile.scala 23:34:@193.4]
  wire [31:0] _GEN_21; // @[RegFile.scala 23:50:@194.4]
  wire  _T_328; // @[RegFile.scala 23:21:@197.4]
  wire  _T_329; // @[RegFile.scala 23:34:@198.4]
  wire [31:0] _GEN_22; // @[RegFile.scala 23:50:@199.4]
  wire  _T_331; // @[RegFile.scala 23:21:@202.4]
  wire  _T_332; // @[RegFile.scala 23:34:@203.4]
  wire [31:0] _GEN_23; // @[RegFile.scala 23:50:@204.4]
  wire  _T_334; // @[RegFile.scala 23:21:@207.4]
  wire  _T_335; // @[RegFile.scala 23:34:@208.4]
  wire [31:0] _GEN_24; // @[RegFile.scala 23:50:@209.4]
  wire  _T_337; // @[RegFile.scala 23:21:@212.4]
  wire  _T_338; // @[RegFile.scala 23:34:@213.4]
  wire [31:0] _GEN_25; // @[RegFile.scala 23:50:@214.4]
  wire  _T_340; // @[RegFile.scala 23:21:@217.4]
  wire  _T_341; // @[RegFile.scala 23:34:@218.4]
  wire [31:0] _GEN_26; // @[RegFile.scala 23:50:@219.4]
  wire  _T_343; // @[RegFile.scala 23:21:@222.4]
  wire  _T_344; // @[RegFile.scala 23:34:@223.4]
  wire [31:0] _GEN_27; // @[RegFile.scala 23:50:@224.4]
  wire  _T_346; // @[RegFile.scala 23:21:@227.4]
  wire  _T_347; // @[RegFile.scala 23:34:@228.4]
  wire [31:0] _GEN_28; // @[RegFile.scala 23:50:@229.4]
  wire  _T_349; // @[RegFile.scala 23:21:@232.4]
  wire  _T_350; // @[RegFile.scala 23:34:@233.4]
  wire [31:0] _GEN_29; // @[RegFile.scala 23:50:@234.4]
  wire  _T_352; // @[RegFile.scala 23:21:@237.4]
  wire  _T_353; // @[RegFile.scala 23:34:@238.4]
  wire [31:0] _GEN_30; // @[RegFile.scala 23:50:@239.4]
  wire  _T_355; // @[RegFile.scala 23:21:@242.4]
  wire  _T_356; // @[RegFile.scala 23:34:@243.4]
  wire [31:0] _GEN_31; // @[RegFile.scala 23:50:@244.4]
  wire  raZero; // @[RegFile.scala 33:27:@247.4]
  wire  rbZero; // @[RegFile.scala 34:27:@248.4]
  wire  rcZero; // @[RegFile.scala 35:27:@249.4]
  wire [31:0] _GEN_33; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_34; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_35; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_36; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_37; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_38; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_39; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_40; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_41; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_42; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_43; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_44; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_45; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_46; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_47; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_48; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_49; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_50; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_51; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_52; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_53; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_54; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_55; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_56; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_57; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_58; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_59; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_60; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_61; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_62; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_63; // @[RegFile.scala 36:19:@250.4]
  wire [31:0] _GEN_65; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_66; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_67; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_68; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_69; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_70; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_71; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_72; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_73; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_74; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_75; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_76; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_77; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_78; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_79; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_80; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_81; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_82; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_83; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_84; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_85; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_86; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_87; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_88; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_89; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_90; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_91; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_92; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_93; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_94; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_95; // @[RegFile.scala 37:19:@252.4]
  wire [31:0] _GEN_97; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_98; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_99; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_100; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_101; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_102; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_103; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_104; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_105; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_106; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_107; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_108; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_109; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_110; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_111; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_112; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_113; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_114; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_115; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_116; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_117; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_118; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_119; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_120; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_121; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_122; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_123; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_124; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_125; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_126; // @[RegFile.scala 38:19:@254.4]
  wire [31:0] _GEN_127; // @[RegFile.scala 38:19:@254.4]
  assign _T_262 = io_wa == 5'h0; // @[RegFile.scala 23:21:@87.4]
  assign _T_263 = _T_262 & io_RegWrite; // @[RegFile.scala 23:34:@88.4]
  assign _GEN_0 = _T_263 ? io_wd : regs_0; // @[RegFile.scala 23:50:@89.4]
  assign _T_265 = io_wa == 5'h1; // @[RegFile.scala 23:21:@92.4]
  assign _T_266 = _T_265 & io_RegWrite; // @[RegFile.scala 23:34:@93.4]
  assign _GEN_1 = _T_266 ? io_wd : regs_1; // @[RegFile.scala 23:50:@94.4]
  assign _T_268 = io_wa == 5'h2; // @[RegFile.scala 23:21:@97.4]
  assign _T_269 = _T_268 & io_RegWrite; // @[RegFile.scala 23:34:@98.4]
  assign _GEN_2 = _T_269 ? io_wd : regs_2; // @[RegFile.scala 23:50:@99.4]
  assign _T_271 = io_wa == 5'h3; // @[RegFile.scala 23:21:@102.4]
  assign _T_272 = _T_271 & io_RegWrite; // @[RegFile.scala 23:34:@103.4]
  assign _GEN_3 = _T_272 ? io_wd : regs_3; // @[RegFile.scala 23:50:@104.4]
  assign _T_274 = io_wa == 5'h4; // @[RegFile.scala 23:21:@107.4]
  assign _T_275 = _T_274 & io_RegWrite; // @[RegFile.scala 23:34:@108.4]
  assign _GEN_4 = _T_275 ? io_wd : regs_4; // @[RegFile.scala 23:50:@109.4]
  assign _T_277 = io_wa == 5'h5; // @[RegFile.scala 23:21:@112.4]
  assign _T_278 = _T_277 & io_RegWrite; // @[RegFile.scala 23:34:@113.4]
  assign _GEN_5 = _T_278 ? io_wd : regs_5; // @[RegFile.scala 23:50:@114.4]
  assign _T_280 = io_wa == 5'h6; // @[RegFile.scala 23:21:@117.4]
  assign _T_281 = _T_280 & io_RegWrite; // @[RegFile.scala 23:34:@118.4]
  assign _GEN_6 = _T_281 ? io_wd : regs_6; // @[RegFile.scala 23:50:@119.4]
  assign _T_283 = io_wa == 5'h7; // @[RegFile.scala 23:21:@122.4]
  assign _T_284 = _T_283 & io_RegWrite; // @[RegFile.scala 23:34:@123.4]
  assign _GEN_7 = _T_284 ? io_wd : regs_7; // @[RegFile.scala 23:50:@124.4]
  assign _T_286 = io_wa == 5'h8; // @[RegFile.scala 23:21:@127.4]
  assign _T_287 = _T_286 & io_RegWrite; // @[RegFile.scala 23:34:@128.4]
  assign _GEN_8 = _T_287 ? io_wd : regs_8; // @[RegFile.scala 23:50:@129.4]
  assign _T_289 = io_wa == 5'h9; // @[RegFile.scala 23:21:@132.4]
  assign _T_290 = _T_289 & io_RegWrite; // @[RegFile.scala 23:34:@133.4]
  assign _GEN_9 = _T_290 ? io_wd : regs_9; // @[RegFile.scala 23:50:@134.4]
  assign _T_292 = io_wa == 5'ha; // @[RegFile.scala 23:21:@137.4]
  assign _T_293 = _T_292 & io_RegWrite; // @[RegFile.scala 23:34:@138.4]
  assign _GEN_10 = _T_293 ? io_wd : regs_10; // @[RegFile.scala 23:50:@139.4]
  assign _T_295 = io_wa == 5'hb; // @[RegFile.scala 23:21:@142.4]
  assign _T_296 = _T_295 & io_RegWrite; // @[RegFile.scala 23:34:@143.4]
  assign _GEN_11 = _T_296 ? io_wd : regs_11; // @[RegFile.scala 23:50:@144.4]
  assign _T_298 = io_wa == 5'hc; // @[RegFile.scala 23:21:@147.4]
  assign _T_299 = _T_298 & io_RegWrite; // @[RegFile.scala 23:34:@148.4]
  assign _GEN_12 = _T_299 ? io_wd : regs_12; // @[RegFile.scala 23:50:@149.4]
  assign _T_301 = io_wa == 5'hd; // @[RegFile.scala 23:21:@152.4]
  assign _T_302 = _T_301 & io_RegWrite; // @[RegFile.scala 23:34:@153.4]
  assign _GEN_13 = _T_302 ? io_wd : regs_13; // @[RegFile.scala 23:50:@154.4]
  assign _T_304 = io_wa == 5'he; // @[RegFile.scala 23:21:@157.4]
  assign _T_305 = _T_304 & io_RegWrite; // @[RegFile.scala 23:34:@158.4]
  assign _GEN_14 = _T_305 ? io_wd : regs_14; // @[RegFile.scala 23:50:@159.4]
  assign _T_307 = io_wa == 5'hf; // @[RegFile.scala 23:21:@162.4]
  assign _T_308 = _T_307 & io_RegWrite; // @[RegFile.scala 23:34:@163.4]
  assign _GEN_15 = _T_308 ? io_wd : regs_15; // @[RegFile.scala 23:50:@164.4]
  assign _T_310 = io_wa == 5'h10; // @[RegFile.scala 23:21:@167.4]
  assign _T_311 = _T_310 & io_RegWrite; // @[RegFile.scala 23:34:@168.4]
  assign _GEN_16 = _T_311 ? io_wd : regs_16; // @[RegFile.scala 23:50:@169.4]
  assign _T_313 = io_wa == 5'h11; // @[RegFile.scala 23:21:@172.4]
  assign _T_314 = _T_313 & io_RegWrite; // @[RegFile.scala 23:34:@173.4]
  assign _GEN_17 = _T_314 ? io_wd : regs_17; // @[RegFile.scala 23:50:@174.4]
  assign _T_316 = io_wa == 5'h12; // @[RegFile.scala 23:21:@177.4]
  assign _T_317 = _T_316 & io_RegWrite; // @[RegFile.scala 23:34:@178.4]
  assign _GEN_18 = _T_317 ? io_wd : regs_18; // @[RegFile.scala 23:50:@179.4]
  assign _T_319 = io_wa == 5'h13; // @[RegFile.scala 23:21:@182.4]
  assign _T_320 = _T_319 & io_RegWrite; // @[RegFile.scala 23:34:@183.4]
  assign _GEN_19 = _T_320 ? io_wd : regs_19; // @[RegFile.scala 23:50:@184.4]
  assign _T_322 = io_wa == 5'h14; // @[RegFile.scala 23:21:@187.4]
  assign _T_323 = _T_322 & io_RegWrite; // @[RegFile.scala 23:34:@188.4]
  assign _GEN_20 = _T_323 ? io_wd : regs_20; // @[RegFile.scala 23:50:@189.4]
  assign _T_325 = io_wa == 5'h15; // @[RegFile.scala 23:21:@192.4]
  assign _T_326 = _T_325 & io_RegWrite; // @[RegFile.scala 23:34:@193.4]
  assign _GEN_21 = _T_326 ? io_wd : regs_21; // @[RegFile.scala 23:50:@194.4]
  assign _T_328 = io_wa == 5'h16; // @[RegFile.scala 23:21:@197.4]
  assign _T_329 = _T_328 & io_RegWrite; // @[RegFile.scala 23:34:@198.4]
  assign _GEN_22 = _T_329 ? io_wd : regs_22; // @[RegFile.scala 23:50:@199.4]
  assign _T_331 = io_wa == 5'h17; // @[RegFile.scala 23:21:@202.4]
  assign _T_332 = _T_331 & io_RegWrite; // @[RegFile.scala 23:34:@203.4]
  assign _GEN_23 = _T_332 ? io_wd : regs_23; // @[RegFile.scala 23:50:@204.4]
  assign _T_334 = io_wa == 5'h18; // @[RegFile.scala 23:21:@207.4]
  assign _T_335 = _T_334 & io_RegWrite; // @[RegFile.scala 23:34:@208.4]
  assign _GEN_24 = _T_335 ? io_wd : regs_24; // @[RegFile.scala 23:50:@209.4]
  assign _T_337 = io_wa == 5'h19; // @[RegFile.scala 23:21:@212.4]
  assign _T_338 = _T_337 & io_RegWrite; // @[RegFile.scala 23:34:@213.4]
  assign _GEN_25 = _T_338 ? io_wd : regs_25; // @[RegFile.scala 23:50:@214.4]
  assign _T_340 = io_wa == 5'h1a; // @[RegFile.scala 23:21:@217.4]
  assign _T_341 = _T_340 & io_RegWrite; // @[RegFile.scala 23:34:@218.4]
  assign _GEN_26 = _T_341 ? io_wd : regs_26; // @[RegFile.scala 23:50:@219.4]
  assign _T_343 = io_wa == 5'h1b; // @[RegFile.scala 23:21:@222.4]
  assign _T_344 = _T_343 & io_RegWrite; // @[RegFile.scala 23:34:@223.4]
  assign _GEN_27 = _T_344 ? io_wd : regs_27; // @[RegFile.scala 23:50:@224.4]
  assign _T_346 = io_wa == 5'h1c; // @[RegFile.scala 23:21:@227.4]
  assign _T_347 = _T_346 & io_RegWrite; // @[RegFile.scala 23:34:@228.4]
  assign _GEN_28 = _T_347 ? io_wd : regs_28; // @[RegFile.scala 23:50:@229.4]
  assign _T_349 = io_wa == 5'h1d; // @[RegFile.scala 23:21:@232.4]
  assign _T_350 = _T_349 & io_RegWrite; // @[RegFile.scala 23:34:@233.4]
  assign _GEN_29 = _T_350 ? io_wd : regs_29; // @[RegFile.scala 23:50:@234.4]
  assign _T_352 = io_wa == 5'h1e; // @[RegFile.scala 23:21:@237.4]
  assign _T_353 = _T_352 & io_RegWrite; // @[RegFile.scala 23:34:@238.4]
  assign _GEN_30 = _T_353 ? io_wd : regs_30; // @[RegFile.scala 23:50:@239.4]
  assign _T_355 = io_wa == 5'h1f; // @[RegFile.scala 23:21:@242.4]
  assign _T_356 = _T_355 & io_RegWrite; // @[RegFile.scala 23:34:@243.4]
  assign _GEN_31 = _T_356 ? io_wd : regs_31; // @[RegFile.scala 23:50:@244.4]
  assign raZero = io_ra_a == 5'h0; // @[RegFile.scala 33:27:@247.4]
  assign rbZero = io_ra_b == 5'h0; // @[RegFile.scala 34:27:@248.4]
  assign rcZero = io_ra_c == 5'h0; // @[RegFile.scala 35:27:@249.4]
  assign _GEN_33 = 5'h1 == io_ra_a ? regs_1 : regs_0; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_34 = 5'h2 == io_ra_a ? regs_2 : _GEN_33; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_35 = 5'h3 == io_ra_a ? regs_3 : _GEN_34; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_36 = 5'h4 == io_ra_a ? regs_4 : _GEN_35; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_37 = 5'h5 == io_ra_a ? regs_5 : _GEN_36; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_38 = 5'h6 == io_ra_a ? regs_6 : _GEN_37; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_39 = 5'h7 == io_ra_a ? regs_7 : _GEN_38; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_40 = 5'h8 == io_ra_a ? regs_8 : _GEN_39; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_41 = 5'h9 == io_ra_a ? regs_9 : _GEN_40; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_42 = 5'ha == io_ra_a ? regs_10 : _GEN_41; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_43 = 5'hb == io_ra_a ? regs_11 : _GEN_42; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_44 = 5'hc == io_ra_a ? regs_12 : _GEN_43; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_45 = 5'hd == io_ra_a ? regs_13 : _GEN_44; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_46 = 5'he == io_ra_a ? regs_14 : _GEN_45; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_47 = 5'hf == io_ra_a ? regs_15 : _GEN_46; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_48 = 5'h10 == io_ra_a ? regs_16 : _GEN_47; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_49 = 5'h11 == io_ra_a ? regs_17 : _GEN_48; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_50 = 5'h12 == io_ra_a ? regs_18 : _GEN_49; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_51 = 5'h13 == io_ra_a ? regs_19 : _GEN_50; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_52 = 5'h14 == io_ra_a ? regs_20 : _GEN_51; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_53 = 5'h15 == io_ra_a ? regs_21 : _GEN_52; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_54 = 5'h16 == io_ra_a ? regs_22 : _GEN_53; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_55 = 5'h17 == io_ra_a ? regs_23 : _GEN_54; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_56 = 5'h18 == io_ra_a ? regs_24 : _GEN_55; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_57 = 5'h19 == io_ra_a ? regs_25 : _GEN_56; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_58 = 5'h1a == io_ra_a ? regs_26 : _GEN_57; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_59 = 5'h1b == io_ra_a ? regs_27 : _GEN_58; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_60 = 5'h1c == io_ra_a ? regs_28 : _GEN_59; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_61 = 5'h1d == io_ra_a ? regs_29 : _GEN_60; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_62 = 5'h1e == io_ra_a ? regs_30 : _GEN_61; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_63 = 5'h1f == io_ra_a ? regs_31 : _GEN_62; // @[RegFile.scala 36:19:@250.4]
  assign _GEN_65 = 5'h1 == io_ra_b ? regs_1 : regs_0; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_66 = 5'h2 == io_ra_b ? regs_2 : _GEN_65; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_67 = 5'h3 == io_ra_b ? regs_3 : _GEN_66; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_68 = 5'h4 == io_ra_b ? regs_4 : _GEN_67; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_69 = 5'h5 == io_ra_b ? regs_5 : _GEN_68; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_70 = 5'h6 == io_ra_b ? regs_6 : _GEN_69; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_71 = 5'h7 == io_ra_b ? regs_7 : _GEN_70; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_72 = 5'h8 == io_ra_b ? regs_8 : _GEN_71; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_73 = 5'h9 == io_ra_b ? regs_9 : _GEN_72; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_74 = 5'ha == io_ra_b ? regs_10 : _GEN_73; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_75 = 5'hb == io_ra_b ? regs_11 : _GEN_74; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_76 = 5'hc == io_ra_b ? regs_12 : _GEN_75; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_77 = 5'hd == io_ra_b ? regs_13 : _GEN_76; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_78 = 5'he == io_ra_b ? regs_14 : _GEN_77; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_79 = 5'hf == io_ra_b ? regs_15 : _GEN_78; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_80 = 5'h10 == io_ra_b ? regs_16 : _GEN_79; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_81 = 5'h11 == io_ra_b ? regs_17 : _GEN_80; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_82 = 5'h12 == io_ra_b ? regs_18 : _GEN_81; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_83 = 5'h13 == io_ra_b ? regs_19 : _GEN_82; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_84 = 5'h14 == io_ra_b ? regs_20 : _GEN_83; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_85 = 5'h15 == io_ra_b ? regs_21 : _GEN_84; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_86 = 5'h16 == io_ra_b ? regs_22 : _GEN_85; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_87 = 5'h17 == io_ra_b ? regs_23 : _GEN_86; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_88 = 5'h18 == io_ra_b ? regs_24 : _GEN_87; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_89 = 5'h19 == io_ra_b ? regs_25 : _GEN_88; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_90 = 5'h1a == io_ra_b ? regs_26 : _GEN_89; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_91 = 5'h1b == io_ra_b ? regs_27 : _GEN_90; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_92 = 5'h1c == io_ra_b ? regs_28 : _GEN_91; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_93 = 5'h1d == io_ra_b ? regs_29 : _GEN_92; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_94 = 5'h1e == io_ra_b ? regs_30 : _GEN_93; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_95 = 5'h1f == io_ra_b ? regs_31 : _GEN_94; // @[RegFile.scala 37:19:@252.4]
  assign _GEN_97 = 5'h1 == io_ra_c ? regs_1 : regs_0; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_98 = 5'h2 == io_ra_c ? regs_2 : _GEN_97; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_99 = 5'h3 == io_ra_c ? regs_3 : _GEN_98; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_100 = 5'h4 == io_ra_c ? regs_4 : _GEN_99; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_101 = 5'h5 == io_ra_c ? regs_5 : _GEN_100; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_102 = 5'h6 == io_ra_c ? regs_6 : _GEN_101; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_103 = 5'h7 == io_ra_c ? regs_7 : _GEN_102; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_104 = 5'h8 == io_ra_c ? regs_8 : _GEN_103; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_105 = 5'h9 == io_ra_c ? regs_9 : _GEN_104; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_106 = 5'ha == io_ra_c ? regs_10 : _GEN_105; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_107 = 5'hb == io_ra_c ? regs_11 : _GEN_106; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_108 = 5'hc == io_ra_c ? regs_12 : _GEN_107; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_109 = 5'hd == io_ra_c ? regs_13 : _GEN_108; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_110 = 5'he == io_ra_c ? regs_14 : _GEN_109; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_111 = 5'hf == io_ra_c ? regs_15 : _GEN_110; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_112 = 5'h10 == io_ra_c ? regs_16 : _GEN_111; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_113 = 5'h11 == io_ra_c ? regs_17 : _GEN_112; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_114 = 5'h12 == io_ra_c ? regs_18 : _GEN_113; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_115 = 5'h13 == io_ra_c ? regs_19 : _GEN_114; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_116 = 5'h14 == io_ra_c ? regs_20 : _GEN_115; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_117 = 5'h15 == io_ra_c ? regs_21 : _GEN_116; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_118 = 5'h16 == io_ra_c ? regs_22 : _GEN_117; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_119 = 5'h17 == io_ra_c ? regs_23 : _GEN_118; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_120 = 5'h18 == io_ra_c ? regs_24 : _GEN_119; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_121 = 5'h19 == io_ra_c ? regs_25 : _GEN_120; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_122 = 5'h1a == io_ra_c ? regs_26 : _GEN_121; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_123 = 5'h1b == io_ra_c ? regs_27 : _GEN_122; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_124 = 5'h1c == io_ra_c ? regs_28 : _GEN_123; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_125 = 5'h1d == io_ra_c ? regs_29 : _GEN_124; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_126 = 5'h1e == io_ra_c ? regs_30 : _GEN_125; // @[RegFile.scala 38:19:@254.4]
  assign _GEN_127 = 5'h1f == io_ra_c ? regs_31 : _GEN_126; // @[RegFile.scala 38:19:@254.4]
  assign io_rd_a = raZero ? 32'h0 : _GEN_63; // @[RegFile.scala 36:13:@251.4]
  assign io_rd_b = rbZero ? 32'h0 : _GEN_95; // @[RegFile.scala 37:13:@253.4]
  assign io_rd_c = rcZero ? 32'h0 : _GEN_127; // @[RegFile.scala 38:13:@255.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 32'h0;
    end else begin
      if (_T_263) begin
        regs_0 <= io_wd;
      end
    end
    if (reset) begin
      regs_1 <= 32'h0;
    end else begin
      if (_T_266) begin
        regs_1 <= io_wd;
      end
    end
    if (reset) begin
      regs_2 <= 32'h0;
    end else begin
      if (_T_269) begin
        regs_2 <= io_wd;
      end
    end
    if (reset) begin
      regs_3 <= 32'h0;
    end else begin
      if (_T_272) begin
        regs_3 <= io_wd;
      end
    end
    if (reset) begin
      regs_4 <= 32'h0;
    end else begin
      if (_T_275) begin
        regs_4 <= io_wd;
      end
    end
    if (reset) begin
      regs_5 <= 32'h0;
    end else begin
      if (_T_278) begin
        regs_5 <= io_wd;
      end
    end
    if (reset) begin
      regs_6 <= 32'h0;
    end else begin
      if (_T_281) begin
        regs_6 <= io_wd;
      end
    end
    if (reset) begin
      regs_7 <= 32'h0;
    end else begin
      if (_T_284) begin
        regs_7 <= io_wd;
      end
    end
    if (reset) begin
      regs_8 <= 32'h0;
    end else begin
      if (_T_287) begin
        regs_8 <= io_wd;
      end
    end
    if (reset) begin
      regs_9 <= 32'h0;
    end else begin
      if (_T_290) begin
        regs_9 <= io_wd;
      end
    end
    if (reset) begin
      regs_10 <= 32'h0;
    end else begin
      if (_T_293) begin
        regs_10 <= io_wd;
      end
    end
    if (reset) begin
      regs_11 <= 32'h0;
    end else begin
      if (_T_296) begin
        regs_11 <= io_wd;
      end
    end
    if (reset) begin
      regs_12 <= 32'h0;
    end else begin
      if (_T_299) begin
        regs_12 <= io_wd;
      end
    end
    if (reset) begin
      regs_13 <= 32'h0;
    end else begin
      if (_T_302) begin
        regs_13 <= io_wd;
      end
    end
    if (reset) begin
      regs_14 <= 32'h0;
    end else begin
      if (_T_305) begin
        regs_14 <= io_wd;
      end
    end
    if (reset) begin
      regs_15 <= 32'h0;
    end else begin
      if (_T_308) begin
        regs_15 <= io_wd;
      end
    end
    if (reset) begin
      regs_16 <= 32'h0;
    end else begin
      if (_T_311) begin
        regs_16 <= io_wd;
      end
    end
    if (reset) begin
      regs_17 <= 32'h0;
    end else begin
      if (_T_314) begin
        regs_17 <= io_wd;
      end
    end
    if (reset) begin
      regs_18 <= 32'h0;
    end else begin
      if (_T_317) begin
        regs_18 <= io_wd;
      end
    end
    if (reset) begin
      regs_19 <= 32'h0;
    end else begin
      if (_T_320) begin
        regs_19 <= io_wd;
      end
    end
    if (reset) begin
      regs_20 <= 32'h0;
    end else begin
      if (_T_323) begin
        regs_20 <= io_wd;
      end
    end
    if (reset) begin
      regs_21 <= 32'h0;
    end else begin
      if (_T_326) begin
        regs_21 <= io_wd;
      end
    end
    if (reset) begin
      regs_22 <= 32'h0;
    end else begin
      if (_T_329) begin
        regs_22 <= io_wd;
      end
    end
    if (reset) begin
      regs_23 <= 32'h0;
    end else begin
      if (_T_332) begin
        regs_23 <= io_wd;
      end
    end
    if (reset) begin
      regs_24 <= 32'h0;
    end else begin
      if (_T_335) begin
        regs_24 <= io_wd;
      end
    end
    if (reset) begin
      regs_25 <= 32'h0;
    end else begin
      if (_T_338) begin
        regs_25 <= io_wd;
      end
    end
    if (reset) begin
      regs_26 <= 32'h0;
    end else begin
      if (_T_341) begin
        regs_26 <= io_wd;
      end
    end
    if (reset) begin
      regs_27 <= 32'h0;
    end else begin
      if (_T_344) begin
        regs_27 <= io_wd;
      end
    end
    if (reset) begin
      regs_28 <= 32'h0;
    end else begin
      if (_T_347) begin
        regs_28 <= io_wd;
      end
    end
    if (reset) begin
      regs_29 <= 32'h0;
    end else begin
      if (_T_350) begin
        regs_29 <= io_wd;
      end
    end
    if (reset) begin
      regs_30 <= 32'h0;
    end else begin
      if (_T_353) begin
        regs_30 <= io_wd;
      end
    end
    if (reset) begin
      regs_31 <= 32'h0;
    end else begin
      if (_T_356) begin
        regs_31 <= io_wd;
      end
    end
  end
endmodule
module Datapath( // @[:@257.2]
  input         clock, // @[:@258.4]
  input         reset, // @[:@259.4]
  output [31:0] io_ctrl_Inst, // @[:@260.4]
  input         io_ctrl_IRWrite, // @[:@260.4]
  input  [1:0]  io_ctrl_RegDst, // @[:@260.4]
  input         io_ctrl_RegWrite, // @[:@260.4]
  input  [1:0]  io_ctrl_ALUSrcA, // @[:@260.4]
  input  [2:0]  io_ctrl_ALUSrcB, // @[:@260.4]
  input  [3:0]  io_ctrl_ALUOp, // @[:@260.4]
  input  [1:0]  io_ctrl_PCSource, // @[:@260.4]
  input         io_ctrl_PCWriteBEQ, // @[:@260.4]
  input         io_ctrl_PCWriteBNE, // @[:@260.4]
  input         io_ctrl_PCWrite, // @[:@260.4]
  input         io_ctrl_IorD, // @[:@260.4]
  input         io_ctrl_MemWrite, // @[:@260.4]
  input  [1:0]  io_ctrl_MemtoReg, // @[:@260.4]
  input  [31:0] io_mem_mem_rdata, // @[:@260.4]
  output [31:0] io_mem_mem_addr, // @[:@260.4]
  output [31:0] io_mem_mem_wdata, // @[:@260.4]
  output        io_mem_mem_wen, // @[:@260.4]
  output [31:0] io_mem_mem_addr2, // @[:@260.4]
  input  [31:0] io_mem_mem_rdata2, // @[:@260.4]
  output [31:0] io_debug_pc, // @[:@260.4]
  input  [4:0]  io_debug_ra_c, // @[:@260.4]
  output [31:0] io_debug_rd_c, // @[:@260.4]
  input  [31:0] io_debug_mr_a, // @[:@260.4]
  output [31:0] io_debug_mr_d // @[:@260.4]
);
  wire [31:0] alu_io_A; // @[Datapath.scala 26:21:@262.4]
  wire [31:0] alu_io_B; // @[Datapath.scala 26:21:@262.4]
  wire [3:0] alu_io_opcode; // @[Datapath.scala 26:21:@262.4]
  wire [31:0] alu_io_out; // @[Datapath.scala 26:21:@262.4]
  wire  alu_io_flagZero; // @[Datapath.scala 26:21:@262.4]
  wire  regFile_clock; // @[Datapath.scala 27:25:@265.4]
  wire  regFile_reset; // @[Datapath.scala 27:25:@265.4]
  wire [4:0] regFile_io_ra_a; // @[Datapath.scala 27:25:@265.4]
  wire [4:0] regFile_io_ra_b; // @[Datapath.scala 27:25:@265.4]
  wire [4:0] regFile_io_wa; // @[Datapath.scala 27:25:@265.4]
  wire [31:0] regFile_io_wd; // @[Datapath.scala 27:25:@265.4]
  wire [31:0] regFile_io_rd_a; // @[Datapath.scala 27:25:@265.4]
  wire [31:0] regFile_io_rd_b; // @[Datapath.scala 27:25:@265.4]
  wire  regFile_io_RegWrite; // @[Datapath.scala 27:25:@265.4]
  wire [4:0] regFile_io_ra_c; // @[Datapath.scala 27:25:@265.4]
  wire [31:0] regFile_io_rd_c; // @[Datapath.scala 27:25:@265.4]
  reg [31:0] ir; // @[Datapath.scala 32:21:@268.4]
  reg [31:0] _RAND_0;
  wire [31:0] _GEN_0; // @[Datapath.scala 33:28:@269.4]
  reg [31:0] mdr; // @[Datapath.scala 39:22:@273.4]
  reg [31:0] _RAND_1;
  reg [31:0] aluout; // @[Datapath.scala 42:25:@275.4]
  reg [31:0] _RAND_2;
  reg [31:0] pc; // @[Datapath.scala 45:21:@277.4]
  reg [31:0] _RAND_3;
  wire  _T_69; // @[Datapath.scala 46:32:@278.4]
  wire  _T_71; // @[Datapath.scala 47:36:@279.4]
  wire  _T_72; // @[Datapath.scala 47:32:@280.4]
  wire  _T_73; // @[Datapath.scala 46:55:@281.4]
  wire  _T_74; // @[Datapath.scala 47:55:@282.4]
  wire [3:0] _T_80; // @[Datapath.scala 52:40:@284.6]
  wire [25:0] _T_81; // @[Datapath.scala 52:52:@285.6]
  wire [27:0] _GEN_2; // @[Datapath.scala 52:59:@286.6]
  wire [27:0] _T_82; // @[Datapath.scala 52:59:@286.6]
  wire [31:0] _T_83; // @[Cat.scala 30:58:@287.6]
  wire  _T_84; // @[Mux.scala 46:19:@288.6]
  wire [31:0] _T_85; // @[Mux.scala 46:16:@289.6]
  wire  _T_86; // @[Mux.scala 46:19:@290.6]
  wire [31:0] _T_87; // @[Mux.scala 46:16:@291.6]
  wire  _T_88; // @[Mux.scala 46:19:@292.6]
  wire [31:0] _T_89; // @[Mux.scala 46:16:@293.6]
  wire  _T_90; // @[Mux.scala 46:19:@294.6]
  wire [31:0] _T_91; // @[Mux.scala 46:16:@295.6]
  wire [31:0] _GEN_1; // @[Datapath.scala 48:31:@283.4]
  wire [4:0] _T_93; // @[Datapath.scala 59:26:@300.4]
  wire [4:0] _T_99; // @[Datapath.scala 63:33:@303.4]
  wire  _T_101; // @[Mux.scala 46:19:@304.4]
  wire [4:0] _T_102; // @[Mux.scala 46:16:@305.4]
  wire  _T_103; // @[Mux.scala 46:19:@306.4]
  wire [4:0] _T_104; // @[Mux.scala 46:16:@307.4]
  wire  _T_105; // @[Mux.scala 46:19:@308.4]
  wire [15:0] _T_112; // @[Datapath.scala 70:45:@311.4]
  wire [31:0] _T_114; // @[Cat.scala 30:58:@312.4]
  wire  _T_115; // @[Mux.scala 46:19:@313.4]
  wire [31:0] _T_116; // @[Mux.scala 46:16:@314.4]
  wire  _T_117; // @[Mux.scala 46:19:@315.4]
  wire [31:0] _T_118; // @[Mux.scala 46:16:@316.4]
  wire  _T_119; // @[Mux.scala 46:19:@317.4]
  wire [31:0] _T_120; // @[Mux.scala 46:16:@318.4]
  wire  _T_121; // @[Mux.scala 46:19:@319.4]
  wire  _T_127; // @[Mux.scala 46:19:@323.4]
  wire [31:0] _T_128; // @[Mux.scala 46:16:@324.4]
  wire  _T_129; // @[Mux.scala 46:19:@325.4]
  wire [31:0] _T_130; // @[Mux.scala 46:16:@326.4]
  wire  _T_131; // @[Mux.scala 46:19:@327.4]
  wire [15:0] _T_144; // @[Datapath.scala 78:16:@332.4]
  wire [31:0] _T_143; // @[Datapath.scala 77:21:@331.4 Datapath.scala 78:11:@333.4]
  wire [31:0] _T_145; // @[Datapath.scala 79:11:@334.4]
  wire [17:0] _GEN_3; // @[Datapath.scala 92:48:@336.4]
  wire [17:0] _T_147; // @[Datapath.scala 92:48:@336.4]
  wire [17:0] _T_150; // @[Datapath.scala 78:16:@338.4]
  wire [31:0] _T_149; // @[Datapath.scala 77:21:@337.4 Datapath.scala 78:11:@339.4]
  wire [31:0] _T_151; // @[Datapath.scala 79:11:@340.4]
  wire [4:0] _T_153; // @[Datapath.scala 94:32:@342.4]
  wire  _T_154; // @[Mux.scala 46:19:@343.4]
  wire [4:0] _T_155; // @[Mux.scala 46:16:@344.4]
  wire  _T_156; // @[Mux.scala 46:19:@345.4]
  wire [15:0] _T_157; // @[Mux.scala 46:16:@346.4]
  wire  _T_158; // @[Mux.scala 46:19:@347.4]
  wire [31:0] _T_159; // @[Mux.scala 46:16:@348.4]
  wire  _T_160; // @[Mux.scala 46:19:@349.4]
  wire [31:0] _T_161; // @[Mux.scala 46:16:@350.4]
  wire  _T_162; // @[Mux.scala 46:19:@351.4]
  wire [31:0] _T_163; // @[Mux.scala 46:16:@352.4]
  wire  _T_164; // @[Mux.scala 46:19:@353.4]
  ALU alu ( // @[Datapath.scala 26:21:@262.4]
    .io_A(alu_io_A),
    .io_B(alu_io_B),
    .io_opcode(alu_io_opcode),
    .io_out(alu_io_out),
    .io_flagZero(alu_io_flagZero)
  );
  RegFile regFile ( // @[Datapath.scala 27:25:@265.4]
    .clock(regFile_clock),
    .reset(regFile_reset),
    .io_ra_a(regFile_io_ra_a),
    .io_ra_b(regFile_io_ra_b),
    .io_wa(regFile_io_wa),
    .io_wd(regFile_io_wd),
    .io_rd_a(regFile_io_rd_a),
    .io_rd_b(regFile_io_rd_b),
    .io_RegWrite(regFile_io_RegWrite),
    .io_ra_c(regFile_io_ra_c),
    .io_rd_c(regFile_io_rd_c)
  );
  assign _GEN_0 = io_ctrl_IRWrite ? io_mem_mem_rdata : ir; // @[Datapath.scala 33:28:@269.4]
  assign _T_69 = io_ctrl_PCWriteBEQ & alu_io_flagZero; // @[Datapath.scala 46:32:@278.4]
  assign _T_71 = alu_io_flagZero == 1'h0; // @[Datapath.scala 47:36:@279.4]
  assign _T_72 = io_ctrl_PCWriteBNE & _T_71; // @[Datapath.scala 47:32:@280.4]
  assign _T_73 = _T_69 | _T_72; // @[Datapath.scala 46:55:@281.4]
  assign _T_74 = _T_73 | io_ctrl_PCWrite; // @[Datapath.scala 47:55:@282.4]
  assign _T_80 = pc[31:28]; // @[Datapath.scala 52:40:@284.6]
  assign _T_81 = ir[25:0]; // @[Datapath.scala 52:52:@285.6]
  assign _GEN_2 = {{2'd0}, _T_81}; // @[Datapath.scala 52:59:@286.6]
  assign _T_82 = _GEN_2 << 2; // @[Datapath.scala 52:59:@286.6]
  assign _T_83 = {_T_80,_T_82}; // @[Cat.scala 30:58:@287.6]
  assign _T_84 = 2'h3 == io_ctrl_PCSource; // @[Mux.scala 46:19:@288.6]
  assign _T_85 = _T_84 ? regFile_io_rd_a : 32'h0; // @[Mux.scala 46:16:@289.6]
  assign _T_86 = 2'h2 == io_ctrl_PCSource; // @[Mux.scala 46:19:@290.6]
  assign _T_87 = _T_86 ? _T_83 : _T_85; // @[Mux.scala 46:16:@291.6]
  assign _T_88 = 2'h1 == io_ctrl_PCSource; // @[Mux.scala 46:19:@292.6]
  assign _T_89 = _T_88 ? aluout : _T_87; // @[Mux.scala 46:16:@293.6]
  assign _T_90 = 2'h0 == io_ctrl_PCSource; // @[Mux.scala 46:19:@294.6]
  assign _T_91 = _T_90 ? alu_io_out : _T_89; // @[Mux.scala 46:16:@295.6]
  assign _GEN_1 = _T_74 ? _T_91 : pc; // @[Datapath.scala 48:31:@283.4]
  assign _T_93 = ir[20:16]; // @[Datapath.scala 59:26:@300.4]
  assign _T_99 = ir[15:11]; // @[Datapath.scala 63:33:@303.4]
  assign _T_101 = 2'h2 == io_ctrl_RegDst; // @[Mux.scala 46:19:@304.4]
  assign _T_102 = _T_101 ? 5'h1f : 5'h0; // @[Mux.scala 46:16:@305.4]
  assign _T_103 = 2'h1 == io_ctrl_RegDst; // @[Mux.scala 46:19:@306.4]
  assign _T_104 = _T_103 ? _T_99 : _T_102; // @[Mux.scala 46:16:@307.4]
  assign _T_105 = 2'h0 == io_ctrl_RegDst; // @[Mux.scala 46:19:@308.4]
  assign _T_112 = ir[15:0]; // @[Datapath.scala 70:45:@311.4]
  assign _T_114 = {_T_112,16'h0}; // @[Cat.scala 30:58:@312.4]
  assign _T_115 = 2'h3 == io_ctrl_MemtoReg; // @[Mux.scala 46:19:@313.4]
  assign _T_116 = _T_115 ? _T_114 : 32'h0; // @[Mux.scala 46:16:@314.4]
  assign _T_117 = 2'h2 == io_ctrl_MemtoReg; // @[Mux.scala 46:19:@315.4]
  assign _T_118 = _T_117 ? pc : _T_116; // @[Mux.scala 46:16:@316.4]
  assign _T_119 = 2'h1 == io_ctrl_MemtoReg; // @[Mux.scala 46:19:@317.4]
  assign _T_120 = _T_119 ? mdr : _T_118; // @[Mux.scala 46:16:@318.4]
  assign _T_121 = 2'h0 == io_ctrl_MemtoReg; // @[Mux.scala 46:19:@319.4]
  assign _T_127 = 2'h2 == io_ctrl_ALUSrcA; // @[Mux.scala 46:19:@323.4]
  assign _T_128 = _T_127 ? regFile_io_rd_b : 32'h0; // @[Mux.scala 46:16:@324.4]
  assign _T_129 = 2'h1 == io_ctrl_ALUSrcA; // @[Mux.scala 46:19:@325.4]
  assign _T_130 = _T_129 ? regFile_io_rd_a : _T_128; // @[Mux.scala 46:16:@326.4]
  assign _T_131 = 2'h0 == io_ctrl_ALUSrcA; // @[Mux.scala 46:19:@327.4]
  assign _T_144 = $signed(_T_112); // @[Datapath.scala 78:16:@332.4]
  assign _T_143 = {{16{_T_144[15]}},_T_144}; // @[Datapath.scala 77:21:@331.4 Datapath.scala 78:11:@333.4]
  assign _T_145 = $unsigned(_T_143); // @[Datapath.scala 79:11:@334.4]
  assign _GEN_3 = {{2'd0}, _T_112}; // @[Datapath.scala 92:48:@336.4]
  assign _T_147 = _GEN_3 << 2; // @[Datapath.scala 92:48:@336.4]
  assign _T_150 = $signed(_T_147); // @[Datapath.scala 78:16:@338.4]
  assign _T_149 = {{14{_T_150[17]}},_T_150}; // @[Datapath.scala 77:21:@337.4 Datapath.scala 78:11:@339.4]
  assign _T_151 = $unsigned(_T_149); // @[Datapath.scala 79:11:@340.4]
  assign _T_153 = ir[10:6]; // @[Datapath.scala 94:32:@342.4]
  assign _T_154 = 3'h5 == io_ctrl_ALUSrcB; // @[Mux.scala 46:19:@343.4]
  assign _T_155 = _T_154 ? _T_153 : 5'h0; // @[Mux.scala 46:16:@344.4]
  assign _T_156 = 3'h4 == io_ctrl_ALUSrcB; // @[Mux.scala 46:19:@345.4]
  assign _T_157 = _T_156 ? _T_112 : {{11'd0}, _T_155}; // @[Mux.scala 46:16:@346.4]
  assign _T_158 = 3'h3 == io_ctrl_ALUSrcB; // @[Mux.scala 46:19:@347.4]
  assign _T_159 = _T_158 ? _T_151 : {{16'd0}, _T_157}; // @[Mux.scala 46:16:@348.4]
  assign _T_160 = 3'h2 == io_ctrl_ALUSrcB; // @[Mux.scala 46:19:@349.4]
  assign _T_161 = _T_160 ? _T_145 : _T_159; // @[Mux.scala 46:16:@350.4]
  assign _T_162 = 3'h1 == io_ctrl_ALUSrcB; // @[Mux.scala 46:19:@351.4]
  assign _T_163 = _T_162 ? 32'h4 : _T_161; // @[Mux.scala 46:16:@352.4]
  assign _T_164 = 3'h0 == io_ctrl_ALUSrcB; // @[Mux.scala 46:19:@353.4]
  assign io_ctrl_Inst = ir; // @[Datapath.scala 36:18:@272.4]
  assign io_mem_mem_addr = io_ctrl_IorD ? aluout : pc; // @[Datapath.scala 101:22:@358.4]
  assign io_mem_mem_wdata = regFile_io_rd_b; // @[Datapath.scala 102:22:@359.4]
  assign io_mem_mem_wen = io_ctrl_MemWrite; // @[Datapath.scala 103:22:@360.4]
  assign io_mem_mem_addr2 = io_debug_mr_a; // @[Datapath.scala 112:22:@367.4]
  assign io_debug_pc = pc; // @[Datapath.scala 109:22:@364.4]
  assign io_debug_rd_c = regFile_io_rd_c; // @[Datapath.scala 111:22:@366.4]
  assign io_debug_mr_d = io_mem_mem_rdata2; // @[Datapath.scala 113:22:@368.4]
  assign alu_io_A = _T_131 ? pc : _T_130; // @[Datapath.scala 83:14:@329.4]
  assign alu_io_B = _T_164 ? regFile_io_rd_b : _T_163; // @[Datapath.scala 88:14:@355.4]
  assign alu_io_opcode = io_ctrl_ALUOp; // @[Datapath.scala 96:19:@356.4]
  assign regFile_clock = clock; // @[:@266.4]
  assign regFile_reset = reset; // @[:@267.4]
  assign regFile_io_ra_a = ir[25:21]; // @[Datapath.scala 58:21:@299.4]
  assign regFile_io_ra_b = ir[20:16]; // @[Datapath.scala 59:21:@301.4]
  assign regFile_io_wa = _T_105 ? _T_93 : _T_104; // @[Datapath.scala 61:21:@310.4]
  assign regFile_io_wd = _T_121 ? aluout : _T_120; // @[Datapath.scala 66:21:@321.4]
  assign regFile_io_RegWrite = io_ctrl_RegWrite; // @[Datapath.scala 74:25:@322.4]
  assign regFile_io_ra_c = io_debug_ra_c; // @[Datapath.scala 110:22:@365.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ir = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mdr = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  aluout = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  pc = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ir <= 32'h20000000;
    end else begin
      if (io_ctrl_IRWrite) begin
        ir <= io_mem_mem_rdata;
      end
    end
    mdr <= io_mem_mem_rdata;
    aluout <= alu_io_out;
    if (reset) begin
      pc <= 32'h0;
    end else begin
      if (_T_74) begin
        if (_T_90) begin
          pc <= alu_io_out;
        end else begin
          if (_T_88) begin
            pc <= aluout;
          end else begin
            if (_T_86) begin
              pc <= _T_83;
            end else begin
              if (_T_84) begin
                pc <= regFile_io_rd_a;
              end else begin
                pc <= 32'h0;
              end
            end
          end
        end
      end
    end
  end
endmodule
module Control( // @[:@370.2]
  input         clock, // @[:@371.4]
  input         reset, // @[:@372.4]
  input  [31:0] io_base_Inst, // @[:@373.4]
  output        io_base_IRWrite, // @[:@373.4]
  output [1:0]  io_base_RegDst, // @[:@373.4]
  output        io_base_RegWrite, // @[:@373.4]
  output [1:0]  io_base_ALUSrcA, // @[:@373.4]
  output [2:0]  io_base_ALUSrcB, // @[:@373.4]
  output [3:0]  io_base_ALUOp, // @[:@373.4]
  output [1:0]  io_base_PCSource, // @[:@373.4]
  output        io_base_PCWriteBEQ, // @[:@373.4]
  output        io_base_PCWriteBNE, // @[:@373.4]
  output        io_base_PCWrite, // @[:@373.4]
  output        io_base_IorD, // @[:@373.4]
  output        io_base_MemWrite, // @[:@373.4]
  output [1:0]  io_base_MemtoReg, // @[:@373.4]
  input         io_SingleStep // @[:@373.4]
);
  wire [31:0] _T_89; // @[Control.scala 156:34:@384.4]
  wire  _T_90; // @[Control.scala 156:34:@385.4]
  wire  _T_94; // @[Control.scala 157:34:@387.4]
  wire  _T_95; // @[Control.scala 156:43:@388.4]
  wire  _T_99; // @[Control.scala 158:34:@390.4]
  wire  _T_100; // @[Control.scala 157:43:@391.4]
  wire  _T_104; // @[Control.scala 159:34:@393.4]
  wire  _T_105; // @[Control.scala 158:43:@394.4]
  wire  _T_109; // @[Control.scala 160:34:@396.4]
  wire  _T_110; // @[Control.scala 159:43:@397.4]
  wire  _T_114; // @[Control.scala 161:34:@399.4]
  wire  _T_115; // @[Control.scala 160:43:@400.4]
  wire  _T_119; // @[Control.scala 162:34:@402.4]
  wire  _T_120; // @[Control.scala 161:43:@403.4]
  wire  _T_124; // @[Control.scala 163:34:@405.4]
  wire  isRType; // @[Control.scala 162:43:@406.4]
  wire [31:0] _T_128; // @[Control.scala 164:31:@408.4]
  wire  _T_129; // @[Control.scala 164:31:@409.4]
  wire  _T_133; // @[Control.scala 165:34:@411.4]
  wire  _T_134; // @[Control.scala 164:41:@412.4]
  wire  _T_138; // @[Control.scala 166:34:@414.4]
  wire  _T_139; // @[Control.scala 165:44:@415.4]
  wire  _T_143; // @[Control.scala 167:34:@417.4]
  wire  _T_144; // @[Control.scala 166:44:@418.4]
  wire  _T_148; // @[Control.scala 168:34:@420.4]
  wire  _T_149; // @[Control.scala 167:44:@421.4]
  wire  _T_153; // @[Control.scala 169:34:@423.4]
  wire  _T_154; // @[Control.scala 168:44:@424.4]
  wire  _T_158; // @[Control.scala 170:34:@426.4]
  wire  isIType; // @[Control.scala 169:45:@427.4]
  wire  _T_163; // @[Control.scala 171:31:@430.4]
  wire  _T_167; // @[Control.scala 171:55:@432.4]
  wire  _T_168; // @[Control.scala 171:38:@433.4]
  wire [31:0] _T_171; // @[Control.scala 171:81:@434.4]
  wire  _T_172; // @[Control.scala 171:81:@435.4]
  wire  isJType; // @[Control.scala 171:64:@436.4]
  wire  isLW; // @[Control.scala 172:30:@439.4]
  wire  isSW; // @[Control.scala 173:30:@442.4]
  wire [31:0] _T_184; // @[Control.scala 174:30:@444.4]
  wire  isLUI; // @[Control.scala 174:30:@445.4]
  wire  isBEQ; // @[Control.scala 175:30:@448.4]
  wire  isBNE; // @[Control.scala 176:30:@451.4]
  wire [31:0] _T_196; // @[Control.scala 177:30:@453.4]
  wire  isSLL; // @[Control.scala 177:30:@454.4]
  reg [4:0] cur_state; // @[Control.scala 198:28:@456.4]
  reg [31:0] _RAND_0;
  wire  _T_212; // @[Conditional.scala 37:30:@471.4]
  wire  _T_218; // @[Control.scala 211:37:@479.6]
  wire [4:0] _T_219; // @[Control.scala 215:32:@482.6]
  wire  _T_220; // @[Conditional.scala 37:30:@486.6]
  wire [4:0] _T_221; // @[Mux.scala 61:16:@491.8]
  wire [4:0] _T_222; // @[Mux.scala 61:16:@492.8]
  wire [4:0] _T_223; // @[Mux.scala 61:16:@493.8]
  wire [4:0] _T_224; // @[Mux.scala 61:16:@494.8]
  wire [4:0] _T_225; // @[Mux.scala 61:16:@495.8]
  wire [4:0] _T_226; // @[Mux.scala 61:16:@496.8]
  wire [4:0] _T_227; // @[Mux.scala 61:16:@497.8]
  wire [4:0] _T_228; // @[Mux.scala 61:16:@498.8]
  wire [4:0] _T_229; // @[Mux.scala 61:16:@499.8]
  wire  _T_230; // @[Conditional.scala 37:30:@503.8]
  wire [4:0] _T_231; // @[Mux.scala 61:16:@508.10]
  wire [4:0] _T_232; // @[Mux.scala 61:16:@509.10]
  wire  _T_233; // @[Conditional.scala 37:30:@513.10]
  wire  _T_236; // @[Conditional.scala 37:30:@523.12]
  wire  _T_239; // @[Conditional.scala 37:30:@533.14]
  wire  _T_242; // @[Conditional.scala 37:30:@540.16]
  wire  _T_245; // @[Conditional.scala 37:30:@547.18]
  wire  _T_247; // @[Conditional.scala 37:30:@555.20]
  wire [3:0] _T_252; // @[Control.scala 117:16:@561.22]
  wire [3:0] _T_257; // @[Control.scala 117:16:@564.22]
  wire [3:0] _T_262; // @[Control.scala 117:16:@567.22]
  wire [3:0] _T_267; // @[Control.scala 117:16:@570.22]
  wire [3:0] _T_272; // @[Control.scala 117:16:@573.22]
  wire [3:0] _T_277; // @[Control.scala 117:16:@576.22]
  wire [3:0] _T_282; // @[Control.scala 117:16:@579.22]
  wire [3:0] _T_287; // @[Control.scala 117:16:@582.22]
  wire  _T_288; // @[Conditional.scala 37:30:@587.22]
  wire  _T_290; // @[Conditional.scala 37:30:@595.24]
  wire  _T_292; // @[Conditional.scala 37:30:@603.26]
  wire [3:0] _T_297; // @[Control.scala 117:16:@609.28]
  wire  _T_298; // @[Conditional.scala 37:30:@614.28]
  wire [2:0] _T_313; // @[Control.scala 117:16:@625.30]
  wire [2:0] _T_318; // @[Control.scala 117:16:@628.30]
  wire [2:0] _T_323; // @[Control.scala 117:16:@631.30]
  wire [2:0] _T_328; // @[Control.scala 117:16:@634.30]
  wire [2:0] _T_333; // @[Control.scala 117:16:@637.30]
  wire [3:0] _T_338; // @[Control.scala 117:16:@641.30]
  wire [3:0] _T_343; // @[Control.scala 117:16:@644.30]
  wire [3:0] _T_348; // @[Control.scala 117:16:@647.30]
  wire [3:0] _T_353; // @[Control.scala 117:16:@650.30]
  wire [3:0] _T_358; // @[Control.scala 117:16:@653.30]
  wire [3:0] _T_363; // @[Control.scala 117:16:@656.30]
  wire [3:0] _T_368; // @[Control.scala 117:16:@659.30]
  wire  _T_369; // @[Conditional.scala 37:30:@664.30]
  wire  _T_371; // @[Conditional.scala 37:30:@672.32]
  wire  _T_372; // @[Conditional.scala 37:30:@683.34]
  wire [1:0] _T_378; // @[Control.scala 117:16:@688.36]
  wire [1:0] _T_383; // @[Control.scala 117:16:@691.36]
  wire [1:0] _T_388; // @[Control.scala 117:16:@694.36]
  wire [1:0] _T_425; // @[Control.scala 117:16:@714.36]
  wire  _T_444; // @[Conditional.scala 37:30:@729.36]
  wire  _T_445; // @[Conditional.scala 37:30:@734.38]
  wire  _T_446; // @[Conditional.scala 37:30:@739.40]
  wire [2:0] _GEN_3; // @[Conditional.scala 39:67:@740.40]
  wire  _GEN_5; // @[Conditional.scala 39:67:@740.40]
  wire [4:0] _GEN_7; // @[Conditional.scala 39:67:@740.40]
  wire [4:0] _GEN_8; // @[Conditional.scala 39:67:@735.38]
  wire  _GEN_9; // @[Conditional.scala 39:67:@735.38]
  wire [2:0] _GEN_12; // @[Conditional.scala 39:67:@735.38]
  wire  _GEN_14; // @[Conditional.scala 39:67:@735.38]
  wire [4:0] _GEN_16; // @[Conditional.scala 39:67:@730.36]
  wire  _GEN_17; // @[Conditional.scala 39:67:@730.36]
  wire [2:0] _GEN_20; // @[Conditional.scala 39:67:@730.36]
  wire  _GEN_22; // @[Conditional.scala 39:67:@730.36]
  wire  _GEN_24; // @[Conditional.scala 39:67:@684.34]
  wire [1:0] _GEN_25; // @[Conditional.scala 39:67:@684.34]
  wire  _GEN_26; // @[Conditional.scala 39:67:@684.34]
  wire [1:0] _GEN_27; // @[Conditional.scala 39:67:@684.34]
  wire [4:0] _GEN_29; // @[Conditional.scala 39:67:@684.34]
  wire  _GEN_30; // @[Conditional.scala 39:67:@684.34]
  wire [2:0] _GEN_33; // @[Conditional.scala 39:67:@684.34]
  wire [1:0] _GEN_35; // @[Conditional.scala 39:67:@673.32]
  wire [2:0] _GEN_36; // @[Conditional.scala 39:67:@673.32]
  wire [3:0] _GEN_37; // @[Conditional.scala 39:67:@673.32]
  wire  _GEN_38; // @[Conditional.scala 39:67:@673.32]
  wire  _GEN_39; // @[Conditional.scala 39:67:@673.32]
  wire [1:0] _GEN_40; // @[Conditional.scala 39:67:@673.32]
  wire [4:0] _GEN_41; // @[Conditional.scala 39:67:@673.32]
  wire  _GEN_42; // @[Conditional.scala 39:67:@673.32]
  wire  _GEN_43; // @[Conditional.scala 39:67:@673.32]
  wire [1:0] _GEN_44; // @[Conditional.scala 39:67:@673.32]
  wire  _GEN_46; // @[Conditional.scala 39:67:@673.32]
  wire [1:0] _GEN_48; // @[Conditional.scala 39:67:@665.30]
  wire  _GEN_49; // @[Conditional.scala 39:67:@665.30]
  wire [4:0] _GEN_51; // @[Conditional.scala 39:67:@665.30]
  wire [1:0] _GEN_52; // @[Conditional.scala 39:67:@665.30]
  wire [2:0] _GEN_53; // @[Conditional.scala 39:67:@665.30]
  wire [3:0] _GEN_54; // @[Conditional.scala 39:67:@665.30]
  wire  _GEN_55; // @[Conditional.scala 39:67:@665.30]
  wire  _GEN_56; // @[Conditional.scala 39:67:@665.30]
  wire [1:0] _GEN_57; // @[Conditional.scala 39:67:@665.30]
  wire  _GEN_58; // @[Conditional.scala 39:67:@665.30]
  wire  _GEN_59; // @[Conditional.scala 39:67:@665.30]
  wire [1:0] _GEN_61; // @[Conditional.scala 39:67:@615.28]
  wire [2:0] _GEN_62; // @[Conditional.scala 39:67:@615.28]
  wire [3:0] _GEN_63; // @[Conditional.scala 39:67:@615.28]
  wire [4:0] _GEN_64; // @[Conditional.scala 39:67:@615.28]
  wire [1:0] _GEN_65; // @[Conditional.scala 39:67:@615.28]
  wire  _GEN_66; // @[Conditional.scala 39:67:@615.28]
  wire  _GEN_68; // @[Conditional.scala 39:67:@615.28]
  wire  _GEN_69; // @[Conditional.scala 39:67:@615.28]
  wire [1:0] _GEN_70; // @[Conditional.scala 39:67:@615.28]
  wire  _GEN_71; // @[Conditional.scala 39:67:@615.28]
  wire  _GEN_72; // @[Conditional.scala 39:67:@615.28]
  wire [1:0] _GEN_74; // @[Conditional.scala 39:67:@604.26]
  wire [2:0] _GEN_75; // @[Conditional.scala 39:67:@604.26]
  wire [3:0] _GEN_76; // @[Conditional.scala 39:67:@604.26]
  wire [4:0] _GEN_77; // @[Conditional.scala 39:67:@604.26]
  wire [1:0] _GEN_78; // @[Conditional.scala 39:67:@604.26]
  wire  _GEN_79; // @[Conditional.scala 39:67:@604.26]
  wire  _GEN_81; // @[Conditional.scala 39:67:@604.26]
  wire  _GEN_82; // @[Conditional.scala 39:67:@604.26]
  wire [1:0] _GEN_83; // @[Conditional.scala 39:67:@604.26]
  wire  _GEN_84; // @[Conditional.scala 39:67:@604.26]
  wire  _GEN_85; // @[Conditional.scala 39:67:@604.26]
  wire [1:0] _GEN_87; // @[Conditional.scala 39:67:@596.24]
  wire  _GEN_88; // @[Conditional.scala 39:67:@596.24]
  wire [1:0] _GEN_89; // @[Conditional.scala 39:67:@596.24]
  wire [4:0] _GEN_90; // @[Conditional.scala 39:67:@596.24]
  wire [1:0] _GEN_91; // @[Conditional.scala 39:67:@596.24]
  wire [2:0] _GEN_92; // @[Conditional.scala 39:67:@596.24]
  wire [3:0] _GEN_93; // @[Conditional.scala 39:67:@596.24]
  wire  _GEN_94; // @[Conditional.scala 39:67:@596.24]
  wire  _GEN_95; // @[Conditional.scala 39:67:@596.24]
  wire [1:0] _GEN_96; // @[Conditional.scala 39:67:@596.24]
  wire  _GEN_97; // @[Conditional.scala 39:67:@596.24]
  wire  _GEN_98; // @[Conditional.scala 39:67:@596.24]
  wire [1:0] _GEN_100; // @[Conditional.scala 39:67:@588.22]
  wire  _GEN_101; // @[Conditional.scala 39:67:@588.22]
  wire [1:0] _GEN_102; // @[Conditional.scala 39:67:@588.22]
  wire [4:0] _GEN_103; // @[Conditional.scala 39:67:@588.22]
  wire [1:0] _GEN_104; // @[Conditional.scala 39:67:@588.22]
  wire [2:0] _GEN_105; // @[Conditional.scala 39:67:@588.22]
  wire [3:0] _GEN_106; // @[Conditional.scala 39:67:@588.22]
  wire  _GEN_107; // @[Conditional.scala 39:67:@588.22]
  wire  _GEN_108; // @[Conditional.scala 39:67:@588.22]
  wire [1:0] _GEN_109; // @[Conditional.scala 39:67:@588.22]
  wire  _GEN_110; // @[Conditional.scala 39:67:@588.22]
  wire  _GEN_111; // @[Conditional.scala 39:67:@588.22]
  wire [1:0] _GEN_113; // @[Conditional.scala 39:67:@556.20]
  wire [2:0] _GEN_114; // @[Conditional.scala 39:67:@556.20]
  wire [3:0] _GEN_115; // @[Conditional.scala 39:67:@556.20]
  wire [4:0] _GEN_116; // @[Conditional.scala 39:67:@556.20]
  wire [1:0] _GEN_117; // @[Conditional.scala 39:67:@556.20]
  wire  _GEN_118; // @[Conditional.scala 39:67:@556.20]
  wire [1:0] _GEN_119; // @[Conditional.scala 39:67:@556.20]
  wire  _GEN_120; // @[Conditional.scala 39:67:@556.20]
  wire  _GEN_121; // @[Conditional.scala 39:67:@556.20]
  wire [1:0] _GEN_122; // @[Conditional.scala 39:67:@556.20]
  wire  _GEN_123; // @[Conditional.scala 39:67:@556.20]
  wire  _GEN_124; // @[Conditional.scala 39:67:@556.20]
  wire [1:0] _GEN_126; // @[Conditional.scala 39:67:@548.18]
  wire  _GEN_127; // @[Conditional.scala 39:67:@548.18]
  wire [1:0] _GEN_128; // @[Conditional.scala 39:67:@548.18]
  wire [4:0] _GEN_129; // @[Conditional.scala 39:67:@548.18]
  wire [1:0] _GEN_130; // @[Conditional.scala 39:67:@548.18]
  wire [2:0] _GEN_131; // @[Conditional.scala 39:67:@548.18]
  wire [3:0] _GEN_132; // @[Conditional.scala 39:67:@548.18]
  wire  _GEN_133; // @[Conditional.scala 39:67:@548.18]
  wire  _GEN_134; // @[Conditional.scala 39:67:@548.18]
  wire [1:0] _GEN_135; // @[Conditional.scala 39:67:@548.18]
  wire  _GEN_136; // @[Conditional.scala 39:67:@548.18]
  wire  _GEN_137; // @[Conditional.scala 39:67:@548.18]
  wire [4:0] _GEN_141; // @[Conditional.scala 39:67:@541.16]
  wire [1:0] _GEN_142; // @[Conditional.scala 39:67:@541.16]
  wire  _GEN_143; // @[Conditional.scala 39:67:@541.16]
  wire [1:0] _GEN_144; // @[Conditional.scala 39:67:@541.16]
  wire [1:0] _GEN_145; // @[Conditional.scala 39:67:@541.16]
  wire [2:0] _GEN_146; // @[Conditional.scala 39:67:@541.16]
  wire [3:0] _GEN_147; // @[Conditional.scala 39:67:@541.16]
  wire  _GEN_148; // @[Conditional.scala 39:67:@541.16]
  wire  _GEN_149; // @[Conditional.scala 39:67:@541.16]
  wire [1:0] _GEN_150; // @[Conditional.scala 39:67:@541.16]
  wire  _GEN_151; // @[Conditional.scala 39:67:@541.16]
  wire  _GEN_152; // @[Conditional.scala 39:67:@541.16]
  wire  _GEN_154; // @[Conditional.scala 39:67:@534.14]
  wire [4:0] _GEN_155; // @[Conditional.scala 39:67:@534.14]
  wire  _GEN_156; // @[Conditional.scala 39:67:@534.14]
  wire [1:0] _GEN_157; // @[Conditional.scala 39:67:@534.14]
  wire  _GEN_158; // @[Conditional.scala 39:67:@534.14]
  wire [1:0] _GEN_159; // @[Conditional.scala 39:67:@534.14]
  wire [1:0] _GEN_160; // @[Conditional.scala 39:67:@534.14]
  wire [2:0] _GEN_161; // @[Conditional.scala 39:67:@534.14]
  wire [3:0] _GEN_162; // @[Conditional.scala 39:67:@534.14]
  wire  _GEN_163; // @[Conditional.scala 39:67:@534.14]
  wire  _GEN_164; // @[Conditional.scala 39:67:@534.14]
  wire [1:0] _GEN_165; // @[Conditional.scala 39:67:@534.14]
  wire  _GEN_166; // @[Conditional.scala 39:67:@534.14]
  wire  _GEN_167; // @[Conditional.scala 39:67:@534.14]
  wire [1:0] _GEN_168; // @[Conditional.scala 39:67:@524.12]
  wire [2:0] _GEN_169; // @[Conditional.scala 39:67:@524.12]
  wire [3:0] _GEN_170; // @[Conditional.scala 39:67:@524.12]
  wire  _GEN_172; // @[Conditional.scala 39:67:@524.12]
  wire [4:0] _GEN_173; // @[Conditional.scala 39:67:@524.12]
  wire  _GEN_174; // @[Conditional.scala 39:67:@524.12]
  wire [1:0] _GEN_175; // @[Conditional.scala 39:67:@524.12]
  wire  _GEN_176; // @[Conditional.scala 39:67:@524.12]
  wire [1:0] _GEN_177; // @[Conditional.scala 39:67:@524.12]
  wire  _GEN_178; // @[Conditional.scala 39:67:@524.12]
  wire  _GEN_179; // @[Conditional.scala 39:67:@524.12]
  wire [1:0] _GEN_180; // @[Conditional.scala 39:67:@524.12]
  wire  _GEN_181; // @[Conditional.scala 39:67:@524.12]
  wire  _GEN_182; // @[Conditional.scala 39:67:@524.12]
  wire [1:0] _GEN_183; // @[Conditional.scala 39:67:@514.10]
  wire [2:0] _GEN_184; // @[Conditional.scala 39:67:@514.10]
  wire [3:0] _GEN_185; // @[Conditional.scala 39:67:@514.10]
  wire  _GEN_187; // @[Conditional.scala 39:67:@514.10]
  wire [4:0] _GEN_188; // @[Conditional.scala 39:67:@514.10]
  wire  _GEN_189; // @[Conditional.scala 39:67:@514.10]
  wire [1:0] _GEN_190; // @[Conditional.scala 39:67:@514.10]
  wire  _GEN_191; // @[Conditional.scala 39:67:@514.10]
  wire [1:0] _GEN_192; // @[Conditional.scala 39:67:@514.10]
  wire  _GEN_193; // @[Conditional.scala 39:67:@514.10]
  wire  _GEN_194; // @[Conditional.scala 39:67:@514.10]
  wire [1:0] _GEN_195; // @[Conditional.scala 39:67:@514.10]
  wire  _GEN_196; // @[Conditional.scala 39:67:@514.10]
  wire  _GEN_197; // @[Conditional.scala 39:67:@514.10]
  wire [1:0] _GEN_198; // @[Conditional.scala 39:67:@504.8]
  wire [2:0] _GEN_199; // @[Conditional.scala 39:67:@504.8]
  wire [3:0] _GEN_200; // @[Conditional.scala 39:67:@504.8]
  wire [4:0] _GEN_201; // @[Conditional.scala 39:67:@504.8]
  wire  _GEN_203; // @[Conditional.scala 39:67:@504.8]
  wire  _GEN_204; // @[Conditional.scala 39:67:@504.8]
  wire [1:0] _GEN_205; // @[Conditional.scala 39:67:@504.8]
  wire  _GEN_206; // @[Conditional.scala 39:67:@504.8]
  wire [1:0] _GEN_207; // @[Conditional.scala 39:67:@504.8]
  wire  _GEN_208; // @[Conditional.scala 39:67:@504.8]
  wire  _GEN_209; // @[Conditional.scala 39:67:@504.8]
  wire [1:0] _GEN_210; // @[Conditional.scala 39:67:@504.8]
  wire  _GEN_211; // @[Conditional.scala 39:67:@504.8]
  wire  _GEN_212; // @[Conditional.scala 39:67:@504.8]
  wire [1:0] _GEN_213; // @[Conditional.scala 39:67:@487.6]
  wire [2:0] _GEN_214; // @[Conditional.scala 39:67:@487.6]
  wire [3:0] _GEN_215; // @[Conditional.scala 39:67:@487.6]
  wire [4:0] _GEN_216; // @[Conditional.scala 39:67:@487.6]
  wire  _GEN_218; // @[Conditional.scala 39:67:@487.6]
  wire  _GEN_219; // @[Conditional.scala 39:67:@487.6]
  wire [1:0] _GEN_220; // @[Conditional.scala 39:67:@487.6]
  wire  _GEN_221; // @[Conditional.scala 39:67:@487.6]
  wire [1:0] _GEN_222; // @[Conditional.scala 39:67:@487.6]
  wire  _GEN_223; // @[Conditional.scala 39:67:@487.6]
  wire  _GEN_224; // @[Conditional.scala 39:67:@487.6]
  wire [1:0] _GEN_225; // @[Conditional.scala 39:67:@487.6]
  wire  _GEN_226; // @[Conditional.scala 39:67:@487.6]
  wire  _GEN_227; // @[Conditional.scala 39:67:@487.6]
  wire [4:0] _GEN_236; // @[Conditional.scala 40:58:@472.4]
  assign _T_89 = io_base_Inst & 32'hfc0007ff; // @[Control.scala 156:34:@384.4]
  assign _T_90 = 32'h20 == _T_89; // @[Control.scala 156:34:@385.4]
  assign _T_94 = 32'h21 == _T_89; // @[Control.scala 157:34:@387.4]
  assign _T_95 = _T_90 | _T_94; // @[Control.scala 156:43:@388.4]
  assign _T_99 = 32'h24 == _T_89; // @[Control.scala 158:34:@390.4]
  assign _T_100 = _T_95 | _T_99; // @[Control.scala 157:43:@391.4]
  assign _T_104 = 32'h22 == _T_89; // @[Control.scala 159:34:@393.4]
  assign _T_105 = _T_100 | _T_104; // @[Control.scala 158:43:@394.4]
  assign _T_109 = 32'h25 == _T_89; // @[Control.scala 160:34:@396.4]
  assign _T_110 = _T_105 | _T_109; // @[Control.scala 159:43:@397.4]
  assign _T_114 = 32'h27 == _T_89; // @[Control.scala 161:34:@399.4]
  assign _T_115 = _T_110 | _T_114; // @[Control.scala 160:43:@400.4]
  assign _T_119 = 32'h26 == _T_89; // @[Control.scala 162:34:@402.4]
  assign _T_120 = _T_115 | _T_119; // @[Control.scala 161:43:@403.4]
  assign _T_124 = 32'h2a == _T_89; // @[Control.scala 163:34:@405.4]
  assign isRType = _T_120 | _T_124; // @[Control.scala 162:43:@406.4]
  assign _T_128 = io_base_Inst & 32'hfc000000; // @[Control.scala 164:31:@408.4]
  assign _T_129 = 32'h20000000 == _T_128; // @[Control.scala 164:31:@409.4]
  assign _T_133 = 32'h30000000 == _T_128; // @[Control.scala 165:34:@411.4]
  assign _T_134 = _T_129 | _T_133; // @[Control.scala 164:41:@412.4]
  assign _T_138 = 32'h34000000 == _T_128; // @[Control.scala 166:34:@414.4]
  assign _T_139 = _T_134 | _T_138; // @[Control.scala 165:44:@415.4]
  assign _T_143 = 32'h38000000 == _T_128; // @[Control.scala 167:34:@417.4]
  assign _T_144 = _T_139 | _T_143; // @[Control.scala 166:44:@418.4]
  assign _T_148 = 32'h28000000 == _T_128; // @[Control.scala 168:34:@420.4]
  assign _T_149 = _T_144 | _T_148; // @[Control.scala 167:44:@421.4]
  assign _T_153 = 32'h24000000 == _T_128; // @[Control.scala 169:34:@423.4]
  assign _T_154 = _T_149 | _T_153; // @[Control.scala 168:44:@424.4]
  assign _T_158 = 32'h2c000000 == _T_128; // @[Control.scala 170:34:@426.4]
  assign isIType = _T_154 | _T_158; // @[Control.scala 169:45:@427.4]
  assign _T_163 = 32'h8000000 == _T_128; // @[Control.scala 171:31:@430.4]
  assign _T_167 = 32'hc000000 == _T_128; // @[Control.scala 171:55:@432.4]
  assign _T_168 = _T_163 | _T_167; // @[Control.scala 171:38:@433.4]
  assign _T_171 = io_base_Inst & 32'hfc1fffff; // @[Control.scala 171:81:@434.4]
  assign _T_172 = 32'h8 == _T_171; // @[Control.scala 171:81:@435.4]
  assign isJType = _T_168 | _T_172; // @[Control.scala 171:64:@436.4]
  assign isLW = 32'h8c000000 == _T_128; // @[Control.scala 172:30:@439.4]
  assign isSW = 32'hac000000 == _T_128; // @[Control.scala 173:30:@442.4]
  assign _T_184 = io_base_Inst & 32'hffe00000; // @[Control.scala 174:30:@444.4]
  assign isLUI = 32'h3c000000 == _T_184; // @[Control.scala 174:30:@445.4]
  assign isBEQ = 32'h10000000 == _T_128; // @[Control.scala 175:30:@448.4]
  assign isBNE = 32'h14000000 == _T_128; // @[Control.scala 176:30:@451.4]
  assign _T_196 = io_base_Inst & 32'hffe0003f; // @[Control.scala 177:30:@453.4]
  assign isSLL = 32'h0 == _T_196; // @[Control.scala 177:30:@454.4]
  assign _T_212 = 5'h0 == cur_state; // @[Conditional.scala 37:30:@471.4]
  assign _T_218 = io_SingleStep ? 1'h0 : 1'h1; // @[Control.scala 211:37:@479.6]
  assign _T_219 = io_SingleStep ? 5'h12 : 5'h1; // @[Control.scala 215:32:@482.6]
  assign _T_220 = 5'h1 == cur_state; // @[Conditional.scala 37:30:@486.6]
  assign _T_221 = isLUI ? 5'ha : 5'h10; // @[Mux.scala 61:16:@491.8]
  assign _T_222 = isSLL ? 5'hf : _T_221; // @[Mux.scala 61:16:@492.8]
  assign _T_223 = isBNE ? 5'hd : _T_222; // @[Mux.scala 61:16:@493.8]
  assign _T_224 = isBEQ ? 5'hd : _T_223; // @[Mux.scala 61:16:@494.8]
  assign _T_225 = isSW ? 5'h2 : _T_224; // @[Mux.scala 61:16:@495.8]
  assign _T_226 = isLW ? 5'h2 : _T_225; // @[Mux.scala 61:16:@496.8]
  assign _T_227 = isJType ? 5'he : _T_226; // @[Mux.scala 61:16:@497.8]
  assign _T_228 = isIType ? 5'hb : _T_227; // @[Mux.scala 61:16:@498.8]
  assign _T_229 = isRType ? 5'h8 : _T_228; // @[Mux.scala 61:16:@499.8]
  assign _T_230 = 5'h2 == cur_state; // @[Conditional.scala 37:30:@503.8]
  assign _T_231 = isSW ? 5'h6 : 5'h10; // @[Mux.scala 61:16:@508.10]
  assign _T_232 = isLW ? 5'h4 : _T_231; // @[Mux.scala 61:16:@509.10]
  assign _T_233 = 5'h4 == cur_state; // @[Conditional.scala 37:30:@513.10]
  assign _T_236 = 5'h6 == cur_state; // @[Conditional.scala 37:30:@523.12]
  assign _T_239 = 5'h3 == cur_state; // @[Conditional.scala 37:30:@533.14]
  assign _T_242 = 5'h5 == cur_state; // @[Conditional.scala 37:30:@540.16]
  assign _T_245 = 5'h7 == cur_state; // @[Conditional.scala 37:30:@547.18]
  assign _T_247 = 5'h8 == cur_state; // @[Conditional.scala 37:30:@555.20]
  assign _T_252 = _T_124 ? 4'h5 : 4'hf; // @[Control.scala 117:16:@561.22]
  assign _T_257 = _T_119 ? 4'h4 : _T_252; // @[Control.scala 117:16:@564.22]
  assign _T_262 = _T_114 ? 4'hc : _T_257; // @[Control.scala 117:16:@567.22]
  assign _T_267 = _T_109 ? 4'h3 : _T_262; // @[Control.scala 117:16:@570.22]
  assign _T_272 = _T_104 ? 4'h1 : _T_267; // @[Control.scala 117:16:@573.22]
  assign _T_277 = _T_99 ? 4'h2 : _T_272; // @[Control.scala 117:16:@576.22]
  assign _T_282 = _T_94 ? 4'h0 : _T_277; // @[Control.scala 117:16:@579.22]
  assign _T_287 = _T_90 ? 4'h0 : _T_282; // @[Control.scala 117:16:@582.22]
  assign _T_288 = 5'h9 == cur_state; // @[Conditional.scala 37:30:@587.22]
  assign _T_290 = 5'ha == cur_state; // @[Conditional.scala 37:30:@595.24]
  assign _T_292 = 5'hf == cur_state; // @[Conditional.scala 37:30:@603.26]
  assign _T_297 = isSLL ? 4'h6 : 4'hf; // @[Control.scala 117:16:@609.28]
  assign _T_298 = 5'hb == cur_state; // @[Conditional.scala 37:30:@614.28]
  assign _T_313 = _T_143 ? 3'h4 : 3'h2; // @[Control.scala 117:16:@625.30]
  assign _T_318 = _T_138 ? 3'h4 : _T_313; // @[Control.scala 117:16:@628.30]
  assign _T_323 = _T_133 ? 3'h4 : _T_318; // @[Control.scala 117:16:@631.30]
  assign _T_328 = _T_153 ? 3'h2 : _T_323; // @[Control.scala 117:16:@634.30]
  assign _T_333 = _T_129 ? 3'h2 : _T_328; // @[Control.scala 117:16:@637.30]
  assign _T_338 = _T_158 ? 4'h7 : 4'hf; // @[Control.scala 117:16:@641.30]
  assign _T_343 = _T_148 ? 4'h5 : _T_338; // @[Control.scala 117:16:@644.30]
  assign _T_348 = _T_143 ? 4'h4 : _T_343; // @[Control.scala 117:16:@647.30]
  assign _T_353 = _T_138 ? 4'h3 : _T_348; // @[Control.scala 117:16:@650.30]
  assign _T_358 = _T_133 ? 4'h2 : _T_353; // @[Control.scala 117:16:@653.30]
  assign _T_363 = _T_153 ? 4'h0 : _T_358; // @[Control.scala 117:16:@656.30]
  assign _T_368 = _T_129 ? 4'h0 : _T_363; // @[Control.scala 117:16:@659.30]
  assign _T_369 = 5'hc == cur_state; // @[Conditional.scala 37:30:@664.30]
  assign _T_371 = 5'hd == cur_state; // @[Conditional.scala 37:30:@672.32]
  assign _T_372 = 5'he == cur_state; // @[Conditional.scala 37:30:@683.34]
  assign _T_378 = _T_172 ? 2'h3 : 2'h2; // @[Control.scala 117:16:@688.36]
  assign _T_383 = _T_163 ? 2'h2 : _T_378; // @[Control.scala 117:16:@691.36]
  assign _T_388 = _T_167 ? 2'h2 : _T_383; // @[Control.scala 117:16:@694.36]
  assign _T_425 = _T_167 ? 2'h2 : 2'h0; // @[Control.scala 117:16:@714.36]
  assign _T_444 = 5'h10 == cur_state; // @[Conditional.scala 37:30:@729.36]
  assign _T_445 = 5'h11 == cur_state; // @[Conditional.scala 37:30:@734.38]
  assign _T_446 = 5'h12 == cur_state; // @[Conditional.scala 37:30:@739.40]
  assign _GEN_3 = _T_446 ? 3'h1 : 3'h0; // @[Conditional.scala 39:67:@740.40]
  assign _GEN_5 = _T_446 ? _T_218 : 1'h0; // @[Conditional.scala 39:67:@740.40]
  assign _GEN_7 = _T_446 ? _T_219 : cur_state; // @[Conditional.scala 39:67:@740.40]
  assign _GEN_8 = _T_445 ? 5'h0 : _GEN_7; // @[Conditional.scala 39:67:@735.38]
  assign _GEN_9 = _T_445 ? 1'h0 : _T_446; // @[Conditional.scala 39:67:@735.38]
  assign _GEN_12 = _T_445 ? 3'h0 : _GEN_3; // @[Conditional.scala 39:67:@735.38]
  assign _GEN_14 = _T_445 ? 1'h0 : _GEN_5; // @[Conditional.scala 39:67:@735.38]
  assign _GEN_16 = _T_444 ? 5'h10 : _GEN_8; // @[Conditional.scala 39:67:@730.36]
  assign _GEN_17 = _T_444 ? 1'h0 : _GEN_9; // @[Conditional.scala 39:67:@730.36]
  assign _GEN_20 = _T_444 ? 3'h0 : _GEN_12; // @[Conditional.scala 39:67:@730.36]
  assign _GEN_22 = _T_444 ? 1'h0 : _GEN_14; // @[Conditional.scala 39:67:@730.36]
  assign _GEN_24 = _T_372 ? 1'h1 : _GEN_22; // @[Conditional.scala 39:67:@684.34]
  assign _GEN_25 = _T_372 ? _T_388 : 2'h0; // @[Conditional.scala 39:67:@684.34]
  assign _GEN_26 = _T_372 ? _T_167 : 1'h0; // @[Conditional.scala 39:67:@684.34]
  assign _GEN_27 = _T_372 ? _T_425 : 2'h0; // @[Conditional.scala 39:67:@684.34]
  assign _GEN_29 = _T_372 ? 5'h0 : _GEN_16; // @[Conditional.scala 39:67:@684.34]
  assign _GEN_30 = _T_372 ? 1'h0 : _GEN_17; // @[Conditional.scala 39:67:@684.34]
  assign _GEN_33 = _T_372 ? 3'h0 : _GEN_20; // @[Conditional.scala 39:67:@684.34]
  assign _GEN_35 = _T_371 ? 2'h1 : 2'h0; // @[Conditional.scala 39:67:@673.32]
  assign _GEN_36 = _T_371 ? 3'h0 : _GEN_33; // @[Conditional.scala 39:67:@673.32]
  assign _GEN_37 = _T_371 ? 4'h1 : 4'h0; // @[Conditional.scala 39:67:@673.32]
  assign _GEN_38 = _T_371 ? isBEQ : 1'h0; // @[Conditional.scala 39:67:@673.32]
  assign _GEN_39 = _T_371 ? isBNE : 1'h0; // @[Conditional.scala 39:67:@673.32]
  assign _GEN_40 = _T_371 ? 2'h1 : _GEN_25; // @[Conditional.scala 39:67:@673.32]
  assign _GEN_41 = _T_371 ? 5'h0 : _GEN_29; // @[Conditional.scala 39:67:@673.32]
  assign _GEN_42 = _T_371 ? 1'h0 : _GEN_24; // @[Conditional.scala 39:67:@673.32]
  assign _GEN_43 = _T_371 ? 1'h0 : _GEN_26; // @[Conditional.scala 39:67:@673.32]
  assign _GEN_44 = _T_371 ? 2'h0 : _GEN_27; // @[Conditional.scala 39:67:@673.32]
  assign _GEN_46 = _T_371 ? 1'h0 : _GEN_30; // @[Conditional.scala 39:67:@673.32]
  assign _GEN_48 = _T_369 ? 2'h0 : _GEN_44; // @[Conditional.scala 39:67:@665.30]
  assign _GEN_49 = _T_369 ? 1'h1 : _GEN_43; // @[Conditional.scala 39:67:@665.30]
  assign _GEN_51 = _T_369 ? 5'h0 : _GEN_41; // @[Conditional.scala 39:67:@665.30]
  assign _GEN_52 = _T_369 ? 2'h0 : _GEN_35; // @[Conditional.scala 39:67:@665.30]
  assign _GEN_53 = _T_369 ? 3'h0 : _GEN_36; // @[Conditional.scala 39:67:@665.30]
  assign _GEN_54 = _T_369 ? 4'h0 : _GEN_37; // @[Conditional.scala 39:67:@665.30]
  assign _GEN_55 = _T_369 ? 1'h0 : _GEN_38; // @[Conditional.scala 39:67:@665.30]
  assign _GEN_56 = _T_369 ? 1'h0 : _GEN_39; // @[Conditional.scala 39:67:@665.30]
  assign _GEN_57 = _T_369 ? 2'h0 : _GEN_40; // @[Conditional.scala 39:67:@665.30]
  assign _GEN_58 = _T_369 ? 1'h0 : _GEN_42; // @[Conditional.scala 39:67:@665.30]
  assign _GEN_59 = _T_369 ? 1'h0 : _GEN_46; // @[Conditional.scala 39:67:@665.30]
  assign _GEN_61 = _T_298 ? 2'h1 : _GEN_52; // @[Conditional.scala 39:67:@615.28]
  assign _GEN_62 = _T_298 ? _T_333 : _GEN_53; // @[Conditional.scala 39:67:@615.28]
  assign _GEN_63 = _T_298 ? _T_368 : _GEN_54; // @[Conditional.scala 39:67:@615.28]
  assign _GEN_64 = _T_298 ? 5'hc : _GEN_51; // @[Conditional.scala 39:67:@615.28]
  assign _GEN_65 = _T_298 ? 2'h0 : _GEN_48; // @[Conditional.scala 39:67:@615.28]
  assign _GEN_66 = _T_298 ? 1'h0 : _GEN_49; // @[Conditional.scala 39:67:@615.28]
  assign _GEN_68 = _T_298 ? 1'h0 : _GEN_55; // @[Conditional.scala 39:67:@615.28]
  assign _GEN_69 = _T_298 ? 1'h0 : _GEN_56; // @[Conditional.scala 39:67:@615.28]
  assign _GEN_70 = _T_298 ? 2'h0 : _GEN_57; // @[Conditional.scala 39:67:@615.28]
  assign _GEN_71 = _T_298 ? 1'h0 : _GEN_58; // @[Conditional.scala 39:67:@615.28]
  assign _GEN_72 = _T_298 ? 1'h0 : _GEN_59; // @[Conditional.scala 39:67:@615.28]
  assign _GEN_74 = _T_292 ? 2'h2 : _GEN_61; // @[Conditional.scala 39:67:@604.26]
  assign _GEN_75 = _T_292 ? 3'h5 : _GEN_62; // @[Conditional.scala 39:67:@604.26]
  assign _GEN_76 = _T_292 ? _T_297 : _GEN_63; // @[Conditional.scala 39:67:@604.26]
  assign _GEN_77 = _T_292 ? 5'h9 : _GEN_64; // @[Conditional.scala 39:67:@604.26]
  assign _GEN_78 = _T_292 ? 2'h0 : _GEN_65; // @[Conditional.scala 39:67:@604.26]
  assign _GEN_79 = _T_292 ? 1'h0 : _GEN_66; // @[Conditional.scala 39:67:@604.26]
  assign _GEN_81 = _T_292 ? 1'h0 : _GEN_68; // @[Conditional.scala 39:67:@604.26]
  assign _GEN_82 = _T_292 ? 1'h0 : _GEN_69; // @[Conditional.scala 39:67:@604.26]
  assign _GEN_83 = _T_292 ? 2'h0 : _GEN_70; // @[Conditional.scala 39:67:@604.26]
  assign _GEN_84 = _T_292 ? 1'h0 : _GEN_71; // @[Conditional.scala 39:67:@604.26]
  assign _GEN_85 = _T_292 ? 1'h0 : _GEN_72; // @[Conditional.scala 39:67:@604.26]
  assign _GEN_87 = _T_290 ? 2'h0 : _GEN_78; // @[Conditional.scala 39:67:@596.24]
  assign _GEN_88 = _T_290 ? 1'h1 : _GEN_79; // @[Conditional.scala 39:67:@596.24]
  assign _GEN_89 = _T_290 ? 2'h3 : _GEN_78; // @[Conditional.scala 39:67:@596.24]
  assign _GEN_90 = _T_290 ? 5'h0 : _GEN_77; // @[Conditional.scala 39:67:@596.24]
  assign _GEN_91 = _T_290 ? 2'h0 : _GEN_74; // @[Conditional.scala 39:67:@596.24]
  assign _GEN_92 = _T_290 ? 3'h0 : _GEN_75; // @[Conditional.scala 39:67:@596.24]
  assign _GEN_93 = _T_290 ? 4'h0 : _GEN_76; // @[Conditional.scala 39:67:@596.24]
  assign _GEN_94 = _T_290 ? 1'h0 : _GEN_81; // @[Conditional.scala 39:67:@596.24]
  assign _GEN_95 = _T_290 ? 1'h0 : _GEN_82; // @[Conditional.scala 39:67:@596.24]
  assign _GEN_96 = _T_290 ? 2'h0 : _GEN_83; // @[Conditional.scala 39:67:@596.24]
  assign _GEN_97 = _T_290 ? 1'h0 : _GEN_84; // @[Conditional.scala 39:67:@596.24]
  assign _GEN_98 = _T_290 ? 1'h0 : _GEN_85; // @[Conditional.scala 39:67:@596.24]
  assign _GEN_100 = _T_288 ? 2'h1 : _GEN_87; // @[Conditional.scala 39:67:@588.22]
  assign _GEN_101 = _T_288 ? 1'h1 : _GEN_88; // @[Conditional.scala 39:67:@588.22]
  assign _GEN_102 = _T_288 ? 2'h0 : _GEN_89; // @[Conditional.scala 39:67:@588.22]
  assign _GEN_103 = _T_288 ? 5'h0 : _GEN_90; // @[Conditional.scala 39:67:@588.22]
  assign _GEN_104 = _T_288 ? 2'h0 : _GEN_91; // @[Conditional.scala 39:67:@588.22]
  assign _GEN_105 = _T_288 ? 3'h0 : _GEN_92; // @[Conditional.scala 39:67:@588.22]
  assign _GEN_106 = _T_288 ? 4'h0 : _GEN_93; // @[Conditional.scala 39:67:@588.22]
  assign _GEN_107 = _T_288 ? 1'h0 : _GEN_94; // @[Conditional.scala 39:67:@588.22]
  assign _GEN_108 = _T_288 ? 1'h0 : _GEN_95; // @[Conditional.scala 39:67:@588.22]
  assign _GEN_109 = _T_288 ? 2'h0 : _GEN_96; // @[Conditional.scala 39:67:@588.22]
  assign _GEN_110 = _T_288 ? 1'h0 : _GEN_97; // @[Conditional.scala 39:67:@588.22]
  assign _GEN_111 = _T_288 ? 1'h0 : _GEN_98; // @[Conditional.scala 39:67:@588.22]
  assign _GEN_113 = _T_247 ? 2'h1 : _GEN_104; // @[Conditional.scala 39:67:@556.20]
  assign _GEN_114 = _T_247 ? 3'h0 : _GEN_105; // @[Conditional.scala 39:67:@556.20]
  assign _GEN_115 = _T_247 ? _T_287 : _GEN_106; // @[Conditional.scala 39:67:@556.20]
  assign _GEN_116 = _T_247 ? 5'h9 : _GEN_103; // @[Conditional.scala 39:67:@556.20]
  assign _GEN_117 = _T_247 ? 2'h0 : _GEN_100; // @[Conditional.scala 39:67:@556.20]
  assign _GEN_118 = _T_247 ? 1'h0 : _GEN_101; // @[Conditional.scala 39:67:@556.20]
  assign _GEN_119 = _T_247 ? 2'h0 : _GEN_102; // @[Conditional.scala 39:67:@556.20]
  assign _GEN_120 = _T_247 ? 1'h0 : _GEN_107; // @[Conditional.scala 39:67:@556.20]
  assign _GEN_121 = _T_247 ? 1'h0 : _GEN_108; // @[Conditional.scala 39:67:@556.20]
  assign _GEN_122 = _T_247 ? 2'h0 : _GEN_109; // @[Conditional.scala 39:67:@556.20]
  assign _GEN_123 = _T_247 ? 1'h0 : _GEN_110; // @[Conditional.scala 39:67:@556.20]
  assign _GEN_124 = _T_247 ? 1'h0 : _GEN_111; // @[Conditional.scala 39:67:@556.20]
  assign _GEN_126 = _T_245 ? 2'h0 : _GEN_117; // @[Conditional.scala 39:67:@548.18]
  assign _GEN_127 = _T_245 ? 1'h1 : _GEN_118; // @[Conditional.scala 39:67:@548.18]
  assign _GEN_128 = _T_245 ? 2'h1 : _GEN_119; // @[Conditional.scala 39:67:@548.18]
  assign _GEN_129 = _T_245 ? 5'h0 : _GEN_116; // @[Conditional.scala 39:67:@548.18]
  assign _GEN_130 = _T_245 ? 2'h0 : _GEN_113; // @[Conditional.scala 39:67:@548.18]
  assign _GEN_131 = _T_245 ? 3'h0 : _GEN_114; // @[Conditional.scala 39:67:@548.18]
  assign _GEN_132 = _T_245 ? 4'h0 : _GEN_115; // @[Conditional.scala 39:67:@548.18]
  assign _GEN_133 = _T_245 ? 1'h0 : _GEN_120; // @[Conditional.scala 39:67:@548.18]
  assign _GEN_134 = _T_245 ? 1'h0 : _GEN_121; // @[Conditional.scala 39:67:@548.18]
  assign _GEN_135 = _T_245 ? 2'h0 : _GEN_122; // @[Conditional.scala 39:67:@548.18]
  assign _GEN_136 = _T_245 ? 1'h0 : _GEN_123; // @[Conditional.scala 39:67:@548.18]
  assign _GEN_137 = _T_245 ? 1'h0 : _GEN_124; // @[Conditional.scala 39:67:@548.18]
  assign _GEN_141 = _T_242 ? 5'h0 : _GEN_129; // @[Conditional.scala 39:67:@541.16]
  assign _GEN_142 = _T_242 ? 2'h0 : _GEN_126; // @[Conditional.scala 39:67:@541.16]
  assign _GEN_143 = _T_242 ? 1'h0 : _GEN_127; // @[Conditional.scala 39:67:@541.16]
  assign _GEN_144 = _T_242 ? 2'h0 : _GEN_128; // @[Conditional.scala 39:67:@541.16]
  assign _GEN_145 = _T_242 ? 2'h0 : _GEN_130; // @[Conditional.scala 39:67:@541.16]
  assign _GEN_146 = _T_242 ? 3'h0 : _GEN_131; // @[Conditional.scala 39:67:@541.16]
  assign _GEN_147 = _T_242 ? 4'h0 : _GEN_132; // @[Conditional.scala 39:67:@541.16]
  assign _GEN_148 = _T_242 ? 1'h0 : _GEN_133; // @[Conditional.scala 39:67:@541.16]
  assign _GEN_149 = _T_242 ? 1'h0 : _GEN_134; // @[Conditional.scala 39:67:@541.16]
  assign _GEN_150 = _T_242 ? 2'h0 : _GEN_135; // @[Conditional.scala 39:67:@541.16]
  assign _GEN_151 = _T_242 ? 1'h0 : _GEN_136; // @[Conditional.scala 39:67:@541.16]
  assign _GEN_152 = _T_242 ? 1'h0 : _GEN_137; // @[Conditional.scala 39:67:@541.16]
  assign _GEN_154 = _T_239 ? 1'h1 : _T_242; // @[Conditional.scala 39:67:@534.14]
  assign _GEN_155 = _T_239 ? 5'h7 : _GEN_141; // @[Conditional.scala 39:67:@534.14]
  assign _GEN_156 = _T_239 ? 1'h0 : _T_242; // @[Conditional.scala 39:67:@534.14]
  assign _GEN_157 = _T_239 ? 2'h0 : _GEN_142; // @[Conditional.scala 39:67:@534.14]
  assign _GEN_158 = _T_239 ? 1'h0 : _GEN_143; // @[Conditional.scala 39:67:@534.14]
  assign _GEN_159 = _T_239 ? 2'h0 : _GEN_144; // @[Conditional.scala 39:67:@534.14]
  assign _GEN_160 = _T_239 ? 2'h0 : _GEN_145; // @[Conditional.scala 39:67:@534.14]
  assign _GEN_161 = _T_239 ? 3'h0 : _GEN_146; // @[Conditional.scala 39:67:@534.14]
  assign _GEN_162 = _T_239 ? 4'h0 : _GEN_147; // @[Conditional.scala 39:67:@534.14]
  assign _GEN_163 = _T_239 ? 1'h0 : _GEN_148; // @[Conditional.scala 39:67:@534.14]
  assign _GEN_164 = _T_239 ? 1'h0 : _GEN_149; // @[Conditional.scala 39:67:@534.14]
  assign _GEN_165 = _T_239 ? 2'h0 : _GEN_150; // @[Conditional.scala 39:67:@534.14]
  assign _GEN_166 = _T_239 ? 1'h0 : _GEN_151; // @[Conditional.scala 39:67:@534.14]
  assign _GEN_167 = _T_239 ? 1'h0 : _GEN_152; // @[Conditional.scala 39:67:@534.14]
  assign _GEN_168 = _T_236 ? 2'h1 : _GEN_160; // @[Conditional.scala 39:67:@524.12]
  assign _GEN_169 = _T_236 ? 3'h2 : _GEN_161; // @[Conditional.scala 39:67:@524.12]
  assign _GEN_170 = _T_236 ? 4'h0 : _GEN_162; // @[Conditional.scala 39:67:@524.12]
  assign _GEN_172 = _T_236 ? 1'h1 : _GEN_154; // @[Conditional.scala 39:67:@524.12]
  assign _GEN_173 = _T_236 ? 5'h5 : _GEN_155; // @[Conditional.scala 39:67:@524.12]
  assign _GEN_174 = _T_236 ? 1'h0 : _GEN_156; // @[Conditional.scala 39:67:@524.12]
  assign _GEN_175 = _T_236 ? 2'h0 : _GEN_157; // @[Conditional.scala 39:67:@524.12]
  assign _GEN_176 = _T_236 ? 1'h0 : _GEN_158; // @[Conditional.scala 39:67:@524.12]
  assign _GEN_177 = _T_236 ? 2'h0 : _GEN_159; // @[Conditional.scala 39:67:@524.12]
  assign _GEN_178 = _T_236 ? 1'h0 : _GEN_163; // @[Conditional.scala 39:67:@524.12]
  assign _GEN_179 = _T_236 ? 1'h0 : _GEN_164; // @[Conditional.scala 39:67:@524.12]
  assign _GEN_180 = _T_236 ? 2'h0 : _GEN_165; // @[Conditional.scala 39:67:@524.12]
  assign _GEN_181 = _T_236 ? 1'h0 : _GEN_166; // @[Conditional.scala 39:67:@524.12]
  assign _GEN_182 = _T_236 ? 1'h0 : _GEN_167; // @[Conditional.scala 39:67:@524.12]
  assign _GEN_183 = _T_233 ? 2'h1 : _GEN_168; // @[Conditional.scala 39:67:@514.10]
  assign _GEN_184 = _T_233 ? 3'h2 : _GEN_169; // @[Conditional.scala 39:67:@514.10]
  assign _GEN_185 = _T_233 ? 4'h0 : _GEN_170; // @[Conditional.scala 39:67:@514.10]
  assign _GEN_187 = _T_233 ? 1'h1 : _GEN_172; // @[Conditional.scala 39:67:@514.10]
  assign _GEN_188 = _T_233 ? 5'h3 : _GEN_173; // @[Conditional.scala 39:67:@514.10]
  assign _GEN_189 = _T_233 ? 1'h0 : _GEN_174; // @[Conditional.scala 39:67:@514.10]
  assign _GEN_190 = _T_233 ? 2'h0 : _GEN_175; // @[Conditional.scala 39:67:@514.10]
  assign _GEN_191 = _T_233 ? 1'h0 : _GEN_176; // @[Conditional.scala 39:67:@514.10]
  assign _GEN_192 = _T_233 ? 2'h0 : _GEN_177; // @[Conditional.scala 39:67:@514.10]
  assign _GEN_193 = _T_233 ? 1'h0 : _GEN_178; // @[Conditional.scala 39:67:@514.10]
  assign _GEN_194 = _T_233 ? 1'h0 : _GEN_179; // @[Conditional.scala 39:67:@514.10]
  assign _GEN_195 = _T_233 ? 2'h0 : _GEN_180; // @[Conditional.scala 39:67:@514.10]
  assign _GEN_196 = _T_233 ? 1'h0 : _GEN_181; // @[Conditional.scala 39:67:@514.10]
  assign _GEN_197 = _T_233 ? 1'h0 : _GEN_182; // @[Conditional.scala 39:67:@514.10]
  assign _GEN_198 = _T_230 ? 2'h1 : _GEN_183; // @[Conditional.scala 39:67:@504.8]
  assign _GEN_199 = _T_230 ? 3'h2 : _GEN_184; // @[Conditional.scala 39:67:@504.8]
  assign _GEN_200 = _T_230 ? 4'h0 : _GEN_185; // @[Conditional.scala 39:67:@504.8]
  assign _GEN_201 = _T_230 ? _T_232 : _GEN_188; // @[Conditional.scala 39:67:@504.8]
  assign _GEN_203 = _T_230 ? 1'h0 : _GEN_187; // @[Conditional.scala 39:67:@504.8]
  assign _GEN_204 = _T_230 ? 1'h0 : _GEN_189; // @[Conditional.scala 39:67:@504.8]
  assign _GEN_205 = _T_230 ? 2'h0 : _GEN_190; // @[Conditional.scala 39:67:@504.8]
  assign _GEN_206 = _T_230 ? 1'h0 : _GEN_191; // @[Conditional.scala 39:67:@504.8]
  assign _GEN_207 = _T_230 ? 2'h0 : _GEN_192; // @[Conditional.scala 39:67:@504.8]
  assign _GEN_208 = _T_230 ? 1'h0 : _GEN_193; // @[Conditional.scala 39:67:@504.8]
  assign _GEN_209 = _T_230 ? 1'h0 : _GEN_194; // @[Conditional.scala 39:67:@504.8]
  assign _GEN_210 = _T_230 ? 2'h0 : _GEN_195; // @[Conditional.scala 39:67:@504.8]
  assign _GEN_211 = _T_230 ? 1'h0 : _GEN_196; // @[Conditional.scala 39:67:@504.8]
  assign _GEN_212 = _T_230 ? 1'h0 : _GEN_197; // @[Conditional.scala 39:67:@504.8]
  assign _GEN_213 = _T_220 ? 2'h0 : _GEN_198; // @[Conditional.scala 39:67:@487.6]
  assign _GEN_214 = _T_220 ? 3'h3 : _GEN_199; // @[Conditional.scala 39:67:@487.6]
  assign _GEN_215 = _T_220 ? 4'h0 : _GEN_200; // @[Conditional.scala 39:67:@487.6]
  assign _GEN_216 = _T_220 ? _T_229 : _GEN_201; // @[Conditional.scala 39:67:@487.6]
  assign _GEN_218 = _T_220 ? 1'h0 : _GEN_203; // @[Conditional.scala 39:67:@487.6]
  assign _GEN_219 = _T_220 ? 1'h0 : _GEN_204; // @[Conditional.scala 39:67:@487.6]
  assign _GEN_220 = _T_220 ? 2'h0 : _GEN_205; // @[Conditional.scala 39:67:@487.6]
  assign _GEN_221 = _T_220 ? 1'h0 : _GEN_206; // @[Conditional.scala 39:67:@487.6]
  assign _GEN_222 = _T_220 ? 2'h0 : _GEN_207; // @[Conditional.scala 39:67:@487.6]
  assign _GEN_223 = _T_220 ? 1'h0 : _GEN_208; // @[Conditional.scala 39:67:@487.6]
  assign _GEN_224 = _T_220 ? 1'h0 : _GEN_209; // @[Conditional.scala 39:67:@487.6]
  assign _GEN_225 = _T_220 ? 2'h0 : _GEN_210; // @[Conditional.scala 39:67:@487.6]
  assign _GEN_226 = _T_220 ? 1'h0 : _GEN_211; // @[Conditional.scala 39:67:@487.6]
  assign _GEN_227 = _T_220 ? 1'h0 : _GEN_212; // @[Conditional.scala 39:67:@487.6]
  assign _GEN_236 = _T_212 ? _T_219 : _GEN_216; // @[Conditional.scala 40:58:@472.4]
  assign io_base_IRWrite = _T_212 ? 1'h1 : _GEN_227; // @[Control.scala 180:30:@457.4 Control.scala 208:31:@476.6 Control.scala 421:31:@744.42]
  assign io_base_RegDst = _T_212 ? 2'h0 : _GEN_220; // @[Control.scala 181:30:@458.4 Control.scala 283:31:@549.20 Control.scala 308:31:@589.24 Control.scala 315:31:@597.26 Control.scala 357:30:@666.32 Control.scala 390:31:@715.36]
  assign io_base_RegWrite = _T_212 ? 1'h0 : _GEN_221; // @[Control.scala 182:30:@459.4 Control.scala 284:31:@550.20 Control.scala 309:31:@590.24 Control.scala 316:31:@598.26 Control.scala 358:31:@667.32 Control.scala 385:31:@705.36]
  assign io_base_ALUSrcA = _T_212 ? 2'h0 : _GEN_213; // @[Control.scala 183:30:@460.4 Control.scala 206:31:@474.6 Control.scala 219:31:@488.8 Control.scala 237:31:@505.10 Control.scala 247:31:@515.12 Control.scala 258:31:@525.14 Control.scala 291:31:@557.22 Control.scala 322:31:@605.28 Control.scala 333:31:@616.30 Control.scala 365:32:@674.34 Control.scala 419:31:@742.42]
  assign io_base_ALUSrcB = _T_212 ? 3'h1 : _GEN_214; // @[Control.scala 184:30:@461.4 Control.scala 209:31:@477.6 Control.scala 220:31:@489.8 Control.scala 238:31:@506.10 Control.scala 248:31:@516.12 Control.scala 259:31:@526.14 Control.scala 292:31:@558.22 Control.scala 323:31:@606.28 Control.scala 334:31:@638.30 Control.scala 366:32:@675.34 Control.scala 422:31:@745.42]
  assign io_base_ALUOp = _T_212 ? 4'h0 : _GEN_215; // @[Control.scala 185:30:@462.4 Control.scala 210:31:@478.6 Control.scala 221:31:@490.8 Control.scala 239:31:@507.10 Control.scala 249:31:@517.12 Control.scala 260:31:@527.14 Control.scala 293:31:@583.22 Control.scala 324:31:@610.28 Control.scala 343:31:@660.30 Control.scala 367:32:@676.34 Control.scala 423:31:@746.42]
  assign io_base_PCSource = _T_212 ? 2'h0 : _GEN_225; // @[Control.scala 186:30:@463.4 Control.scala 212:31:@481.6 Control.scala 370:32:@679.34 Control.scala 379:31:@695.36 Control.scala 426:31:@749.42]
  assign io_base_PCWriteBEQ = _T_212 ? 1'h0 : _GEN_223; // @[Control.scala 187:30:@464.4 Control.scala 368:32:@677.34]
  assign io_base_PCWriteBNE = _T_212 ? 1'h0 : _GEN_224; // @[Control.scala 188:30:@465.4 Control.scala 369:32:@678.34]
  assign io_base_PCWrite = _T_212 ? _T_218 : _GEN_226; // @[Control.scala 189:30:@466.4 Control.scala 211:31:@480.6 Control.scala 377:31:@685.36 Control.scala 425:31:@748.42]
  assign io_base_IorD = _T_212 ? 1'h0 : _GEN_218; // @[Control.scala 190:30:@467.4 Control.scala 207:31:@475.6 Control.scala 252:31:@519.12 Control.scala 263:31:@529.14 Control.scala 270:31:@536.16 Control.scala 277:31:@543.18 Control.scala 420:31:@743.42]
  assign io_base_MemWrite = _T_212 ? 1'h0 : _GEN_219; // @[Control.scala 192:30:@469.4 Control.scala 276:31:@542.18]
  assign io_base_MemtoReg = _T_212 ? 2'h0 : _GEN_222; // @[Control.scala 193:30:@470.4 Control.scala 285:31:@551.20 Control.scala 310:31:@591.24 Control.scala 317:31:@599.26 Control.scala 359:31:@668.32 Control.scala 396:31:@725.36]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cur_state = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cur_state <= 5'h11;
    end else begin
      if (_T_212) begin
        if (io_SingleStep) begin
          cur_state <= 5'h12;
        end else begin
          cur_state <= 5'h1;
        end
      end else begin
        if (_T_220) begin
          if (isRType) begin
            cur_state <= 5'h8;
          end else begin
            if (isIType) begin
              cur_state <= 5'hb;
            end else begin
              if (isJType) begin
                cur_state <= 5'he;
              end else begin
                if (isLW) begin
                  cur_state <= 5'h2;
                end else begin
                  if (isSW) begin
                    cur_state <= 5'h2;
                  end else begin
                    if (isBEQ) begin
                      cur_state <= 5'hd;
                    end else begin
                      if (isBNE) begin
                        cur_state <= 5'hd;
                      end else begin
                        if (isSLL) begin
                          cur_state <= 5'hf;
                        end else begin
                          if (isLUI) begin
                            cur_state <= 5'ha;
                          end else begin
                            cur_state <= 5'h10;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_230) begin
            if (isLW) begin
              cur_state <= 5'h4;
            end else begin
              if (isSW) begin
                cur_state <= 5'h6;
              end else begin
                cur_state <= 5'h10;
              end
            end
          end else begin
            if (_T_233) begin
              cur_state <= 5'h3;
            end else begin
              if (_T_236) begin
                cur_state <= 5'h5;
              end else begin
                if (_T_239) begin
                  cur_state <= 5'h7;
                end else begin
                  if (_T_242) begin
                    cur_state <= 5'h0;
                  end else begin
                    if (_T_245) begin
                      cur_state <= 5'h0;
                    end else begin
                      if (_T_247) begin
                        cur_state <= 5'h9;
                      end else begin
                        if (_T_288) begin
                          cur_state <= 5'h0;
                        end else begin
                          if (_T_290) begin
                            cur_state <= 5'h0;
                          end else begin
                            if (_T_292) begin
                              cur_state <= 5'h9;
                            end else begin
                              if (_T_298) begin
                                cur_state <= 5'hc;
                              end else begin
                                if (_T_369) begin
                                  cur_state <= 5'h0;
                                end else begin
                                  if (_T_371) begin
                                    cur_state <= 5'h0;
                                  end else begin
                                    if (_T_372) begin
                                      cur_state <= 5'h0;
                                    end else begin
                                      if (_T_444) begin
                                        cur_state <= 5'h10;
                                      end else begin
                                        if (_T_445) begin
                                          cur_state <= 5'h0;
                                        end else begin
                                          if (_T_446) begin
                                            if (io_SingleStep) begin
                                              cur_state <= 5'h12;
                                            end else begin
                                              cur_state <= 5'h1;
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module CPU( // @[:@762.2]
  input         clock, // @[:@763.4]
  input         reset, // @[:@764.4]
  output [31:0] io_debug_pc, // @[:@765.4]
  input  [4:0]  io_debug_ra_c, // @[:@765.4]
  output [31:0] io_debug_rd_c, // @[:@765.4]
  input  [31:0] io_debug_mr_a, // @[:@765.4]
  output [31:0] io_debug_mr_d, // @[:@765.4]
  input  [31:0] io_mem_port_mem_rdata, // @[:@765.4]
  output [31:0] io_mem_port_mem_addr, // @[:@765.4]
  output [31:0] io_mem_port_mem_wdata, // @[:@765.4]
  output        io_mem_port_mem_wen, // @[:@765.4]
  output [31:0] io_mem_port_mem_addr2, // @[:@765.4]
  input  [31:0] io_mem_port_mem_rdata2, // @[:@765.4]
  input         io_single // @[:@765.4]
);
  wire  datapath_clock; // @[CPU.scala 15:26:@767.4]
  wire  datapath_reset; // @[CPU.scala 15:26:@767.4]
  wire [31:0] datapath_io_ctrl_Inst; // @[CPU.scala 15:26:@767.4]
  wire  datapath_io_ctrl_IRWrite; // @[CPU.scala 15:26:@767.4]
  wire [1:0] datapath_io_ctrl_RegDst; // @[CPU.scala 15:26:@767.4]
  wire  datapath_io_ctrl_RegWrite; // @[CPU.scala 15:26:@767.4]
  wire [1:0] datapath_io_ctrl_ALUSrcA; // @[CPU.scala 15:26:@767.4]
  wire [2:0] datapath_io_ctrl_ALUSrcB; // @[CPU.scala 15:26:@767.4]
  wire [3:0] datapath_io_ctrl_ALUOp; // @[CPU.scala 15:26:@767.4]
  wire [1:0] datapath_io_ctrl_PCSource; // @[CPU.scala 15:26:@767.4]
  wire  datapath_io_ctrl_PCWriteBEQ; // @[CPU.scala 15:26:@767.4]
  wire  datapath_io_ctrl_PCWriteBNE; // @[CPU.scala 15:26:@767.4]
  wire  datapath_io_ctrl_PCWrite; // @[CPU.scala 15:26:@767.4]
  wire  datapath_io_ctrl_IorD; // @[CPU.scala 15:26:@767.4]
  wire  datapath_io_ctrl_MemWrite; // @[CPU.scala 15:26:@767.4]
  wire [1:0] datapath_io_ctrl_MemtoReg; // @[CPU.scala 15:26:@767.4]
  wire [31:0] datapath_io_mem_mem_rdata; // @[CPU.scala 15:26:@767.4]
  wire [31:0] datapath_io_mem_mem_addr; // @[CPU.scala 15:26:@767.4]
  wire [31:0] datapath_io_mem_mem_wdata; // @[CPU.scala 15:26:@767.4]
  wire  datapath_io_mem_mem_wen; // @[CPU.scala 15:26:@767.4]
  wire [31:0] datapath_io_mem_mem_addr2; // @[CPU.scala 15:26:@767.4]
  wire [31:0] datapath_io_mem_mem_rdata2; // @[CPU.scala 15:26:@767.4]
  wire [31:0] datapath_io_debug_pc; // @[CPU.scala 15:26:@767.4]
  wire [4:0] datapath_io_debug_ra_c; // @[CPU.scala 15:26:@767.4]
  wire [31:0] datapath_io_debug_rd_c; // @[CPU.scala 15:26:@767.4]
  wire [31:0] datapath_io_debug_mr_a; // @[CPU.scala 15:26:@767.4]
  wire [31:0] datapath_io_debug_mr_d; // @[CPU.scala 15:26:@767.4]
  wire  ctrl_clock; // @[CPU.scala 18:22:@778.4]
  wire  ctrl_reset; // @[CPU.scala 18:22:@778.4]
  wire [31:0] ctrl_io_base_Inst; // @[CPU.scala 18:22:@778.4]
  wire  ctrl_io_base_IRWrite; // @[CPU.scala 18:22:@778.4]
  wire [1:0] ctrl_io_base_RegDst; // @[CPU.scala 18:22:@778.4]
  wire  ctrl_io_base_RegWrite; // @[CPU.scala 18:22:@778.4]
  wire [1:0] ctrl_io_base_ALUSrcA; // @[CPU.scala 18:22:@778.4]
  wire [2:0] ctrl_io_base_ALUSrcB; // @[CPU.scala 18:22:@778.4]
  wire [3:0] ctrl_io_base_ALUOp; // @[CPU.scala 18:22:@778.4]
  wire [1:0] ctrl_io_base_PCSource; // @[CPU.scala 18:22:@778.4]
  wire  ctrl_io_base_PCWriteBEQ; // @[CPU.scala 18:22:@778.4]
  wire  ctrl_io_base_PCWriteBNE; // @[CPU.scala 18:22:@778.4]
  wire  ctrl_io_base_PCWrite; // @[CPU.scala 18:22:@778.4]
  wire  ctrl_io_base_IorD; // @[CPU.scala 18:22:@778.4]
  wire  ctrl_io_base_MemWrite; // @[CPU.scala 18:22:@778.4]
  wire [1:0] ctrl_io_base_MemtoReg; // @[CPU.scala 18:22:@778.4]
  wire  ctrl_io_SingleStep; // @[CPU.scala 18:22:@778.4]
  Datapath datapath ( // @[CPU.scala 15:26:@767.4]
    .clock(datapath_clock),
    .reset(datapath_reset),
    .io_ctrl_Inst(datapath_io_ctrl_Inst),
    .io_ctrl_IRWrite(datapath_io_ctrl_IRWrite),
    .io_ctrl_RegDst(datapath_io_ctrl_RegDst),
    .io_ctrl_RegWrite(datapath_io_ctrl_RegWrite),
    .io_ctrl_ALUSrcA(datapath_io_ctrl_ALUSrcA),
    .io_ctrl_ALUSrcB(datapath_io_ctrl_ALUSrcB),
    .io_ctrl_ALUOp(datapath_io_ctrl_ALUOp),
    .io_ctrl_PCSource(datapath_io_ctrl_PCSource),
    .io_ctrl_PCWriteBEQ(datapath_io_ctrl_PCWriteBEQ),
    .io_ctrl_PCWriteBNE(datapath_io_ctrl_PCWriteBNE),
    .io_ctrl_PCWrite(datapath_io_ctrl_PCWrite),
    .io_ctrl_IorD(datapath_io_ctrl_IorD),
    .io_ctrl_MemWrite(datapath_io_ctrl_MemWrite),
    .io_ctrl_MemtoReg(datapath_io_ctrl_MemtoReg),
    .io_mem_mem_rdata(datapath_io_mem_mem_rdata),
    .io_mem_mem_addr(datapath_io_mem_mem_addr),
    .io_mem_mem_wdata(datapath_io_mem_mem_wdata),
    .io_mem_mem_wen(datapath_io_mem_mem_wen),
    .io_mem_mem_addr2(datapath_io_mem_mem_addr2),
    .io_mem_mem_rdata2(datapath_io_mem_mem_rdata2),
    .io_debug_pc(datapath_io_debug_pc),
    .io_debug_ra_c(datapath_io_debug_ra_c),
    .io_debug_rd_c(datapath_io_debug_rd_c),
    .io_debug_mr_a(datapath_io_debug_mr_a),
    .io_debug_mr_d(datapath_io_debug_mr_d)
  );
  Control ctrl ( // @[CPU.scala 18:22:@778.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_base_Inst(ctrl_io_base_Inst),
    .io_base_IRWrite(ctrl_io_base_IRWrite),
    .io_base_RegDst(ctrl_io_base_RegDst),
    .io_base_RegWrite(ctrl_io_base_RegWrite),
    .io_base_ALUSrcA(ctrl_io_base_ALUSrcA),
    .io_base_ALUSrcB(ctrl_io_base_ALUSrcB),
    .io_base_ALUOp(ctrl_io_base_ALUOp),
    .io_base_PCSource(ctrl_io_base_PCSource),
    .io_base_PCWriteBEQ(ctrl_io_base_PCWriteBEQ),
    .io_base_PCWriteBNE(ctrl_io_base_PCWriteBNE),
    .io_base_PCWrite(ctrl_io_base_PCWrite),
    .io_base_IorD(ctrl_io_base_IorD),
    .io_base_MemWrite(ctrl_io_base_MemWrite),
    .io_base_MemtoReg(ctrl_io_base_MemtoReg),
    .io_SingleStep(ctrl_io_SingleStep)
  );
  assign io_debug_pc = datapath_io_debug_pc; // @[CPU.scala 16:14:@774.4]
  assign io_debug_rd_c = datapath_io_debug_rd_c; // @[CPU.scala 16:14:@772.4]
  assign io_debug_mr_d = datapath_io_debug_mr_d; // @[CPU.scala 16:14:@770.4]
  assign io_mem_port_mem_addr = datapath_io_mem_mem_addr; // @[CPU.scala 23:17:@809.4]
  assign io_mem_port_mem_wdata = datapath_io_mem_mem_wdata; // @[CPU.scala 23:17:@808.4]
  assign io_mem_port_mem_wen = datapath_io_mem_mem_wen; // @[CPU.scala 23:17:@807.4]
  assign io_mem_port_mem_addr2 = datapath_io_mem_mem_addr2; // @[CPU.scala 23:17:@806.4]
  assign datapath_clock = clock; // @[:@768.4]
  assign datapath_reset = reset; // @[:@769.4]
  assign datapath_io_ctrl_IRWrite = ctrl_io_base_IRWrite; // @[CPU.scala 19:18:@794.4]
  assign datapath_io_ctrl_RegDst = ctrl_io_base_RegDst; // @[CPU.scala 19:18:@793.4]
  assign datapath_io_ctrl_RegWrite = ctrl_io_base_RegWrite; // @[CPU.scala 19:18:@792.4]
  assign datapath_io_ctrl_ALUSrcA = ctrl_io_base_ALUSrcA; // @[CPU.scala 19:18:@791.4]
  assign datapath_io_ctrl_ALUSrcB = ctrl_io_base_ALUSrcB; // @[CPU.scala 19:18:@790.4]
  assign datapath_io_ctrl_ALUOp = ctrl_io_base_ALUOp; // @[CPU.scala 19:18:@789.4]
  assign datapath_io_ctrl_PCSource = ctrl_io_base_PCSource; // @[CPU.scala 19:18:@788.4]
  assign datapath_io_ctrl_PCWriteBEQ = ctrl_io_base_PCWriteBEQ; // @[CPU.scala 19:18:@787.4]
  assign datapath_io_ctrl_PCWriteBNE = ctrl_io_base_PCWriteBNE; // @[CPU.scala 19:18:@786.4]
  assign datapath_io_ctrl_PCWrite = ctrl_io_base_PCWrite; // @[CPU.scala 19:18:@785.4]
  assign datapath_io_ctrl_IorD = ctrl_io_base_IorD; // @[CPU.scala 19:18:@784.4]
  assign datapath_io_ctrl_MemWrite = ctrl_io_base_MemWrite; // @[CPU.scala 19:18:@782.4]
  assign datapath_io_ctrl_MemtoReg = ctrl_io_base_MemtoReg; // @[CPU.scala 19:18:@781.4]
  assign datapath_io_mem_mem_rdata = io_mem_port_mem_rdata; // @[CPU.scala 23:17:@810.4]
  assign datapath_io_mem_mem_rdata2 = io_mem_port_mem_rdata2; // @[CPU.scala 23:17:@805.4]
  assign datapath_io_debug_ra_c = io_debug_ra_c; // @[CPU.scala 16:14:@773.4]
  assign datapath_io_debug_mr_a = io_debug_mr_a; // @[CPU.scala 16:14:@771.4]
  assign ctrl_clock = clock; // @[:@779.4]
  assign ctrl_reset = reset; // @[:@780.4]
  assign ctrl_io_base_Inst = datapath_io_ctrl_Inst; // @[CPU.scala 19:18:@795.4]
  assign ctrl_io_SingleStep = io_single; // @[CPU.scala 21:24:@804.4]
endmodule
module MMap( // @[:@812.2]
  output [31:0] io_mmap_port_mem_rdata, // @[:@815.4]
  input  [31:0] io_mmap_port_mem_addr, // @[:@815.4]
  input  [31:0] io_mmap_port_mem_wdata, // @[:@815.4]
  input         io_mmap_port_mem_wen, // @[:@815.4]
  input  [31:0] io_mmap_port_mem_addr2, // @[:@815.4]
  output [31:0] io_mmap_port_mem_rdata2, // @[:@815.4]
  input  [31:0] io_mem_port_mem_rdata, // @[:@815.4]
  output [31:0] io_mem_port_mem_addr, // @[:@815.4]
  output [31:0] io_mem_port_mem_wdata, // @[:@815.4]
  output        io_mem_port_mem_wen, // @[:@815.4]
  output [31:0] io_mem_port_mem_addr2, // @[:@815.4]
  input  [31:0] io_mem_port_mem_rdata2, // @[:@815.4]
  input  [31:0] io_uart_port_mem_rdata, // @[:@815.4]
  output [31:0] io_uart_port_mem_wdata, // @[:@815.4]
  output        io_uart_port_mem_wen, // @[:@815.4]
  output [31:0] io_vram_port_mem_addr, // @[:@815.4]
  output [15:0] io_vram_port_mem_wdata, // @[:@815.4]
  output        io_vram_port_mem_wen // @[:@815.4]
);
  wire  addr_in_mem; // @[MMap.scala 46:81:@818.4]
  wire  addr_in_uart; // @[MMap.scala 47:47:@820.4]
  wire  _T_61; // @[MMap.scala 48:47:@821.4]
  wire  _T_63; // @[MMap.scala 48:85:@822.4]
  wire  addr_in_vram; // @[MMap.scala 48:59:@823.4]
  wire [31:0] _T_67; // @[Mux.scala 61:16:@825.4]
  wire [32:0] _T_72; // @[MMap.scala 68:53:@837.4]
  wire [32:0] _T_73; // @[MMap.scala 68:53:@838.4]
  wire [31:0] _T_74; // @[MMap.scala 68:53:@839.4]
  wire [29:0] _T_75; // @[MMap.scala 68:64:@840.4]
  assign addr_in_mem = io_mmap_port_mem_addr < 32'h400; // @[MMap.scala 46:81:@818.4]
  assign addr_in_uart = io_mmap_port_mem_addr == 32'hff00; // @[MMap.scala 47:47:@820.4]
  assign _T_61 = io_mmap_port_mem_addr >= 32'h3000; // @[MMap.scala 48:47:@821.4]
  assign _T_63 = io_mmap_port_mem_addr < 32'h4f41; // @[MMap.scala 48:85:@822.4]
  assign addr_in_vram = _T_61 & _T_63; // @[MMap.scala 48:59:@823.4]
  assign _T_67 = addr_in_uart ? io_uart_port_mem_rdata : 32'h0; // @[Mux.scala 61:16:@825.4]
  assign _T_72 = io_mmap_port_mem_addr - 32'h3000; // @[MMap.scala 68:53:@837.4]
  assign _T_73 = $unsigned(_T_72); // @[MMap.scala 68:53:@838.4]
  assign _T_74 = _T_73[31:0]; // @[MMap.scala 68:53:@839.4]
  assign _T_75 = _T_74[31:2]; // @[MMap.scala 68:64:@840.4]
  assign io_mmap_port_mem_rdata = addr_in_mem ? io_mem_port_mem_rdata : _T_67; // @[MMap.scala 50:28:@827.4]
  assign io_mmap_port_mem_rdata2 = io_mem_port_mem_rdata2; // @[MMap.scala 62:29:@833.4]
  assign io_mem_port_mem_addr = io_mmap_port_mem_addr; // @[MMap.scala 57:27:@828.4]
  assign io_mem_port_mem_wdata = io_mmap_port_mem_wdata; // @[MMap.scala 58:27:@829.4]
  assign io_mem_port_mem_wen = io_mmap_port_mem_wen & addr_in_mem; // @[MMap.scala 59:27:@831.4]
  assign io_mem_port_mem_addr2 = io_mmap_port_mem_addr2; // @[MMap.scala 60:27:@832.4]
  assign io_uart_port_mem_wdata = io_mmap_port_mem_wdata; // @[MMap.scala 65:28:@834.4]
  assign io_uart_port_mem_wen = io_mmap_port_mem_wen & addr_in_uart; // @[MMap.scala 66:28:@836.4]
  assign io_vram_port_mem_addr = {{2'd0}, _T_75}; // @[MMap.scala 68:27:@841.4]
  assign io_vram_port_mem_wdata = io_mmap_port_mem_wdata[15:0]; // @[MMap.scala 69:28:@843.4]
  assign io_vram_port_mem_wen = io_mmap_port_mem_wen & addr_in_vram; // @[MMap.scala 70:28:@845.4]
endmodule
module Mem( // @[:@847.2]
  input         clock, // @[:@848.4]
  input         reset, // @[:@849.4]
  output [31:0] io_mem_rdata, // @[:@850.4]
  input  [31:0] io_mem_addr, // @[:@850.4]
  input  [31:0] io_mem_wdata, // @[:@850.4]
  input         io_mem_wen, // @[:@850.4]
  input  [31:0] io_mem_addr2, // @[:@850.4]
  output [31:0] io_mem_rdata2 // @[:@850.4]
);
  reg [31:0] memory_0; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_0;
  reg [31:0] memory_1; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_1;
  reg [31:0] memory_2; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_2;
  reg [31:0] memory_3; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_3;
  reg [31:0] memory_4; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_4;
  reg [31:0] memory_5; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_5;
  reg [31:0] memory_6; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_6;
  reg [31:0] memory_7; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_7;
  reg [31:0] memory_8; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_8;
  reg [31:0] memory_9; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_9;
  reg [31:0] memory_10; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_10;
  reg [31:0] memory_11; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_11;
  reg [31:0] memory_12; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_12;
  reg [31:0] memory_13; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_13;
  reg [31:0] memory_14; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_14;
  reg [31:0] memory_15; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_15;
  reg [31:0] memory_16; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_16;
  reg [31:0] memory_17; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_17;
  reg [31:0] memory_18; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_18;
  reg [31:0] memory_19; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_19;
  reg [31:0] memory_20; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_20;
  reg [31:0] memory_21; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_21;
  reg [31:0] memory_22; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_22;
  reg [31:0] memory_23; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_23;
  reg [31:0] memory_24; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_24;
  reg [31:0] memory_25; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_25;
  reg [31:0] memory_26; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_26;
  reg [31:0] memory_27; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_27;
  reg [31:0] memory_28; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_28;
  reg [31:0] memory_29; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_29;
  reg [31:0] memory_30; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_30;
  reg [31:0] memory_31; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_31;
  reg [31:0] memory_32; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_32;
  reg [31:0] memory_33; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_33;
  reg [31:0] memory_34; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_34;
  reg [31:0] memory_35; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_35;
  reg [31:0] memory_36; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_36;
  reg [31:0] memory_37; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_37;
  reg [31:0] memory_38; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_38;
  reg [31:0] memory_39; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_39;
  reg [31:0] memory_40; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_40;
  reg [31:0] memory_41; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_41;
  reg [31:0] memory_42; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_42;
  reg [31:0] memory_43; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_43;
  reg [31:0] memory_44; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_44;
  reg [31:0] memory_45; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_45;
  reg [31:0] memory_46; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_46;
  reg [31:0] memory_47; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_47;
  reg [31:0] memory_48; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_48;
  reg [31:0] memory_49; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_49;
  reg [31:0] memory_50; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_50;
  reg [31:0] memory_51; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_51;
  reg [31:0] memory_52; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_52;
  reg [31:0] memory_53; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_53;
  reg [31:0] memory_54; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_54;
  reg [31:0] memory_55; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_55;
  reg [31:0] memory_56; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_56;
  reg [31:0] memory_57; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_57;
  reg [31:0] memory_58; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_58;
  reg [31:0] memory_59; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_59;
  reg [31:0] memory_60; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_60;
  reg [31:0] memory_61; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_61;
  reg [31:0] memory_62; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_62;
  reg [31:0] memory_63; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_63;
  reg [31:0] memory_64; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_64;
  reg [31:0] memory_65; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_65;
  reg [31:0] memory_66; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_66;
  reg [31:0] memory_67; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_67;
  reg [31:0] memory_68; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_68;
  reg [31:0] memory_69; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_69;
  reg [31:0] memory_70; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_70;
  reg [31:0] memory_71; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_71;
  reg [31:0] memory_72; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_72;
  reg [31:0] memory_73; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_73;
  reg [31:0] memory_74; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_74;
  reg [31:0] memory_75; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_75;
  reg [31:0] memory_76; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_76;
  reg [31:0] memory_77; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_77;
  reg [31:0] memory_78; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_78;
  reg [31:0] memory_79; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_79;
  reg [31:0] memory_80; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_80;
  reg [31:0] memory_81; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_81;
  reg [31:0] memory_82; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_82;
  reg [31:0] memory_83; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_83;
  reg [31:0] memory_84; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_84;
  reg [31:0] memory_85; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_85;
  reg [31:0] memory_86; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_86;
  reg [31:0] memory_87; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_87;
  reg [31:0] memory_88; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_88;
  reg [31:0] memory_89; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_89;
  reg [31:0] memory_90; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_90;
  reg [31:0] memory_91; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_91;
  reg [31:0] memory_92; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_92;
  reg [31:0] memory_93; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_93;
  reg [31:0] memory_94; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_94;
  reg [31:0] memory_95; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_95;
  reg [31:0] memory_96; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_96;
  reg [31:0] memory_97; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_97;
  reg [31:0] memory_98; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_98;
  reg [31:0] memory_99; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_99;
  reg [31:0] memory_100; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_100;
  reg [31:0] memory_101; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_101;
  reg [31:0] memory_102; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_102;
  reg [31:0] memory_103; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_103;
  reg [31:0] memory_104; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_104;
  reg [31:0] memory_105; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_105;
  reg [31:0] memory_106; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_106;
  reg [31:0] memory_107; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_107;
  reg [31:0] memory_108; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_108;
  reg [31:0] memory_109; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_109;
  reg [31:0] memory_110; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_110;
  reg [31:0] memory_111; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_111;
  reg [31:0] memory_112; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_112;
  reg [31:0] memory_113; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_113;
  reg [31:0] memory_114; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_114;
  reg [31:0] memory_115; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_115;
  reg [31:0] memory_116; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_116;
  reg [31:0] memory_117; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_117;
  reg [31:0] memory_118; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_118;
  reg [31:0] memory_119; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_119;
  reg [31:0] memory_120; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_120;
  reg [31:0] memory_121; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_121;
  reg [31:0] memory_122; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_122;
  reg [31:0] memory_123; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_123;
  reg [31:0] memory_124; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_124;
  reg [31:0] memory_125; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_125;
  reg [31:0] memory_126; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_126;
  reg [31:0] memory_127; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_127;
  reg [31:0] memory_128; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_128;
  reg [31:0] memory_129; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_129;
  reg [31:0] memory_130; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_130;
  reg [31:0] memory_131; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_131;
  reg [31:0] memory_132; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_132;
  reg [31:0] memory_133; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_133;
  reg [31:0] memory_134; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_134;
  reg [31:0] memory_135; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_135;
  reg [31:0] memory_136; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_136;
  reg [31:0] memory_137; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_137;
  reg [31:0] memory_138; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_138;
  reg [31:0] memory_139; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_139;
  reg [31:0] memory_140; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_140;
  reg [31:0] memory_141; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_141;
  reg [31:0] memory_142; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_142;
  reg [31:0] memory_143; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_143;
  reg [31:0] memory_144; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_144;
  reg [31:0] memory_145; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_145;
  reg [31:0] memory_146; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_146;
  reg [31:0] memory_147; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_147;
  reg [31:0] memory_148; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_148;
  reg [31:0] memory_149; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_149;
  reg [31:0] memory_150; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_150;
  reg [31:0] memory_151; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_151;
  reg [31:0] memory_152; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_152;
  reg [31:0] memory_153; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_153;
  reg [31:0] memory_154; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_154;
  reg [31:0] memory_155; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_155;
  reg [31:0] memory_156; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_156;
  reg [31:0] memory_157; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_157;
  reg [31:0] memory_158; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_158;
  reg [31:0] memory_159; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_159;
  reg [31:0] memory_160; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_160;
  reg [31:0] memory_161; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_161;
  reg [31:0] memory_162; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_162;
  reg [31:0] memory_163; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_163;
  reg [31:0] memory_164; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_164;
  reg [31:0] memory_165; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_165;
  reg [31:0] memory_166; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_166;
  reg [31:0] memory_167; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_167;
  reg [31:0] memory_168; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_168;
  reg [31:0] memory_169; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_169;
  reg [31:0] memory_170; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_170;
  reg [31:0] memory_171; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_171;
  reg [31:0] memory_172; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_172;
  reg [31:0] memory_173; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_173;
  reg [31:0] memory_174; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_174;
  reg [31:0] memory_175; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_175;
  reg [31:0] memory_176; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_176;
  reg [31:0] memory_177; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_177;
  reg [31:0] memory_178; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_178;
  reg [31:0] memory_179; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_179;
  reg [31:0] memory_180; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_180;
  reg [31:0] memory_181; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_181;
  reg [31:0] memory_182; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_182;
  reg [31:0] memory_183; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_183;
  reg [31:0] memory_184; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_184;
  reg [31:0] memory_185; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_185;
  reg [31:0] memory_186; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_186;
  reg [31:0] memory_187; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_187;
  reg [31:0] memory_188; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_188;
  reg [31:0] memory_189; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_189;
  reg [31:0] memory_190; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_190;
  reg [31:0] memory_191; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_191;
  reg [31:0] memory_192; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_192;
  reg [31:0] memory_193; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_193;
  reg [31:0] memory_194; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_194;
  reg [31:0] memory_195; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_195;
  reg [31:0] memory_196; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_196;
  reg [31:0] memory_197; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_197;
  reg [31:0] memory_198; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_198;
  reg [31:0] memory_199; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_199;
  reg [31:0] memory_200; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_200;
  reg [31:0] memory_201; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_201;
  reg [31:0] memory_202; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_202;
  reg [31:0] memory_203; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_203;
  reg [31:0] memory_204; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_204;
  reg [31:0] memory_205; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_205;
  reg [31:0] memory_206; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_206;
  reg [31:0] memory_207; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_207;
  reg [31:0] memory_208; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_208;
  reg [31:0] memory_209; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_209;
  reg [31:0] memory_210; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_210;
  reg [31:0] memory_211; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_211;
  reg [31:0] memory_212; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_212;
  reg [31:0] memory_213; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_213;
  reg [31:0] memory_214; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_214;
  reg [31:0] memory_215; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_215;
  reg [31:0] memory_216; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_216;
  reg [31:0] memory_217; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_217;
  reg [31:0] memory_218; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_218;
  reg [31:0] memory_219; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_219;
  reg [31:0] memory_220; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_220;
  reg [31:0] memory_221; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_221;
  reg [31:0] memory_222; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_222;
  reg [31:0] memory_223; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_223;
  reg [31:0] memory_224; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_224;
  reg [31:0] memory_225; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_225;
  reg [31:0] memory_226; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_226;
  reg [31:0] memory_227; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_227;
  reg [31:0] memory_228; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_228;
  reg [31:0] memory_229; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_229;
  reg [31:0] memory_230; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_230;
  reg [31:0] memory_231; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_231;
  reg [31:0] memory_232; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_232;
  reg [31:0] memory_233; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_233;
  reg [31:0] memory_234; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_234;
  reg [31:0] memory_235; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_235;
  reg [31:0] memory_236; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_236;
  reg [31:0] memory_237; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_237;
  reg [31:0] memory_238; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_238;
  reg [31:0] memory_239; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_239;
  reg [31:0] memory_240; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_240;
  reg [31:0] memory_241; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_241;
  reg [31:0] memory_242; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_242;
  reg [31:0] memory_243; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_243;
  reg [31:0] memory_244; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_244;
  reg [31:0] memory_245; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_245;
  reg [31:0] memory_246; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_246;
  reg [31:0] memory_247; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_247;
  reg [31:0] memory_248; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_248;
  reg [31:0] memory_249; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_249;
  reg [31:0] memory_250; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_250;
  reg [31:0] memory_251; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_251;
  reg [31:0] memory_252; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_252;
  reg [31:0] memory_253; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_253;
  reg [31:0] memory_254; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_254;
  reg [31:0] memory_255; // @[Mem.scala 58:25:@1109.4]
  reg [31:0] _RAND_255;
  wire [29:0] _T_1830; // @[Mem.scala 65:28:@1111.6]
  wire [7:0] _T_1834; // @[:@1112.6]
  wire [31:0] _GEN_0; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_1; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_2; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_3; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_4; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_5; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_6; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_7; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_8; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_9; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_10; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_11; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_12; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_13; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_14; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_15; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_16; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_17; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_18; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_19; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_20; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_21; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_22; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_23; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_24; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_25; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_26; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_27; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_28; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_29; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_30; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_31; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_32; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_33; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_34; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_35; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_36; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_37; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_38; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_39; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_40; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_41; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_42; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_43; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_44; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_45; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_46; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_47; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_48; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_49; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_50; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_51; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_52; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_53; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_54; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_55; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_56; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_57; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_58; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_59; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_60; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_61; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_62; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_63; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_64; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_65; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_66; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_67; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_68; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_69; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_70; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_71; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_72; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_73; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_74; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_75; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_76; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_77; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_78; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_79; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_80; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_81; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_82; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_83; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_84; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_85; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_86; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_87; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_88; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_89; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_90; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_91; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_92; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_93; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_94; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_95; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_96; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_97; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_98; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_99; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_100; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_101; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_102; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_103; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_104; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_105; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_106; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_107; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_108; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_109; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_110; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_111; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_112; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_113; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_114; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_115; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_116; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_117; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_118; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_119; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_120; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_121; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_122; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_123; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_124; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_125; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_126; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_127; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_128; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_129; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_130; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_131; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_132; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_133; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_134; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_135; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_136; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_137; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_138; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_139; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_140; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_141; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_142; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_143; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_144; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_145; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_146; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_147; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_148; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_149; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_150; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_151; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_152; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_153; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_154; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_155; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_156; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_157; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_158; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_159; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_160; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_161; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_162; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_163; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_164; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_165; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_166; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_167; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_168; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_169; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_170; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_171; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_172; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_173; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_174; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_175; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_176; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_177; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_178; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_179; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_180; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_181; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_182; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_183; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_184; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_185; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_186; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_187; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_188; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_189; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_190; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_191; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_192; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_193; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_194; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_195; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_196; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_197; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_198; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_199; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_200; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_201; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_202; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_203; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_204; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_205; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_206; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_207; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_208; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_209; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_210; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_211; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_212; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_213; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_214; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_215; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_216; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_217; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_218; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_219; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_220; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_221; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_222; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_223; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_224; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_225; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_226; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_227; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_228; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_229; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_230; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_231; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_232; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_233; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_234; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_235; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_236; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_237; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_238; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_239; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_240; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_241; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_242; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_243; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_244; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_245; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_246; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_247; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_248; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_249; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_250; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_251; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_252; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_253; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_254; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_255; // @[Mem.scala 65:34:@1113.6]
  wire [31:0] _GEN_256; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_257; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_258; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_259; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_260; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_261; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_262; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_263; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_264; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_265; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_266; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_267; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_268; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_269; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_270; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_271; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_272; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_273; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_274; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_275; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_276; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_277; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_278; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_279; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_280; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_281; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_282; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_283; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_284; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_285; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_286; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_287; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_288; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_289; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_290; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_291; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_292; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_293; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_294; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_295; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_296; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_297; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_298; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_299; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_300; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_301; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_302; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_303; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_304; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_305; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_306; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_307; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_308; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_309; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_310; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_311; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_312; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_313; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_314; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_315; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_316; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_317; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_318; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_319; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_320; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_321; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_322; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_323; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_324; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_325; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_326; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_327; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_328; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_329; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_330; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_331; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_332; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_333; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_334; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_335; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_336; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_337; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_338; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_339; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_340; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_341; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_342; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_343; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_344; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_345; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_346; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_347; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_348; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_349; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_350; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_351; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_352; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_353; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_354; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_355; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_356; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_357; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_358; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_359; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_360; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_361; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_362; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_363; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_364; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_365; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_366; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_367; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_368; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_369; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_370; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_371; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_372; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_373; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_374; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_375; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_376; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_377; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_378; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_379; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_380; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_381; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_382; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_383; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_384; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_385; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_386; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_387; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_388; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_389; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_390; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_391; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_392; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_393; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_394; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_395; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_396; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_397; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_398; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_399; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_400; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_401; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_402; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_403; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_404; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_405; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_406; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_407; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_408; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_409; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_410; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_411; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_412; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_413; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_414; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_415; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_416; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_417; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_418; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_419; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_420; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_421; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_422; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_423; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_424; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_425; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_426; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_427; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_428; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_429; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_430; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_431; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_432; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_433; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_434; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_435; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_436; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_437; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_438; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_439; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_440; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_441; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_442; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_443; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_444; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_445; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_446; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_447; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_448; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_449; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_450; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_451; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_452; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_453; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_454; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_455; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_456; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_457; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_458; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_459; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_460; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_461; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_462; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_463; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_464; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_465; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_466; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_467; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_468; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_469; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_470; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_471; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_472; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_473; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_474; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_475; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_476; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_477; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_478; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_479; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_480; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_481; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_482; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_483; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_484; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_485; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_486; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_487; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_488; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_489; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_490; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_491; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_492; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_493; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_494; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_495; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_496; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_497; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_498; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_499; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_500; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_501; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_502; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_503; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_504; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_505; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_506; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_507; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_508; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_509; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_510; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_511; // @[Mem.scala 64:23:@1110.4]
  wire [31:0] _GEN_513; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_514; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_515; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_516; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_517; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_518; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_519; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_520; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_521; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_522; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_523; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_524; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_525; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_526; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_527; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_528; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_529; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_530; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_531; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_532; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_533; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_534; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_535; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_536; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_537; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_538; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_539; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_540; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_541; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_542; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_543; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_544; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_545; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_546; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_547; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_548; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_549; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_550; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_551; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_552; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_553; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_554; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_555; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_556; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_557; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_558; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_559; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_560; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_561; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_562; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_563; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_564; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_565; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_566; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_567; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_568; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_569; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_570; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_571; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_572; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_573; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_574; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_575; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_576; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_577; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_578; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_579; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_580; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_581; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_582; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_583; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_584; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_585; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_586; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_587; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_588; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_589; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_590; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_591; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_592; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_593; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_594; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_595; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_596; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_597; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_598; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_599; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_600; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_601; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_602; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_603; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_604; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_605; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_606; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_607; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_608; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_609; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_610; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_611; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_612; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_613; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_614; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_615; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_616; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_617; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_618; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_619; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_620; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_621; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_622; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_623; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_624; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_625; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_626; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_627; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_628; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_629; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_630; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_631; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_632; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_633; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_634; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_635; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_636; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_637; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_638; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_639; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_640; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_641; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_642; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_643; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_644; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_645; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_646; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_647; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_648; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_649; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_650; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_651; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_652; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_653; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_654; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_655; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_656; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_657; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_658; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_659; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_660; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_661; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_662; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_663; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_664; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_665; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_666; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_667; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_668; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_669; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_670; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_671; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_672; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_673; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_674; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_675; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_676; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_677; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_678; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_679; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_680; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_681; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_682; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_683; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_684; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_685; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_686; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_687; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_688; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_689; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_690; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_691; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_692; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_693; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_694; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_695; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_696; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_697; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_698; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_699; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_700; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_701; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_702; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_703; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_704; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_705; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_706; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_707; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_708; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_709; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_710; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_711; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_712; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_713; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_714; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_715; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_716; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_717; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_718; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_719; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_720; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_721; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_722; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_723; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_724; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_725; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_726; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_727; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_728; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_729; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_730; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_731; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_732; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_733; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_734; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_735; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_736; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_737; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_738; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_739; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_740; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_741; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_742; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_743; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_744; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_745; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_746; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_747; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_748; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_749; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_750; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_751; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_752; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_753; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_754; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_755; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_756; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_757; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_758; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_759; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_760; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_761; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_762; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_763; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_764; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_765; // @[Mem.scala 69:18:@1117.4]
  wire [31:0] _GEN_766; // @[Mem.scala 69:18:@1117.4]
  wire [29:0] _T_1840; // @[Mem.scala 73:42:@1118.4]
  wire [7:0] _T_1844; // @[:@1119.4]
  wire [31:0] _GEN_769; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_770; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_771; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_772; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_773; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_774; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_775; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_776; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_777; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_778; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_779; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_780; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_781; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_782; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_783; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_784; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_785; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_786; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_787; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_788; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_789; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_790; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_791; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_792; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_793; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_794; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_795; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_796; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_797; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_798; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_799; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_800; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_801; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_802; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_803; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_804; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_805; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_806; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_807; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_808; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_809; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_810; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_811; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_812; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_813; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_814; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_815; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_816; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_817; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_818; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_819; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_820; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_821; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_822; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_823; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_824; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_825; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_826; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_827; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_828; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_829; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_830; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_831; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_832; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_833; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_834; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_835; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_836; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_837; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_838; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_839; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_840; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_841; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_842; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_843; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_844; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_845; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_846; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_847; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_848; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_849; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_850; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_851; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_852; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_853; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_854; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_855; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_856; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_857; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_858; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_859; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_860; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_861; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_862; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_863; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_864; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_865; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_866; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_867; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_868; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_869; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_870; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_871; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_872; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_873; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_874; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_875; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_876; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_877; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_878; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_879; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_880; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_881; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_882; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_883; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_884; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_885; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_886; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_887; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_888; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_889; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_890; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_891; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_892; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_893; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_894; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_895; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_896; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_897; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_898; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_899; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_900; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_901; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_902; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_903; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_904; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_905; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_906; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_907; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_908; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_909; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_910; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_911; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_912; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_913; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_914; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_915; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_916; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_917; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_918; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_919; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_920; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_921; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_922; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_923; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_924; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_925; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_926; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_927; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_928; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_929; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_930; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_931; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_932; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_933; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_934; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_935; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_936; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_937; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_938; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_939; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_940; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_941; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_942; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_943; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_944; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_945; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_946; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_947; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_948; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_949; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_950; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_951; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_952; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_953; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_954; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_955; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_956; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_957; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_958; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_959; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_960; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_961; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_962; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_963; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_964; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_965; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_966; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_967; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_968; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_969; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_970; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_971; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_972; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_973; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_974; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_975; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_976; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_977; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_978; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_979; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_980; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_981; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_982; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_983; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_984; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_985; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_986; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_987; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_988; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_989; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_990; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_991; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_992; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_993; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_994; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_995; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_996; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_997; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_998; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_999; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1000; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1001; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1002; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1003; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1004; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1005; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1006; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1007; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1008; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1009; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1010; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1011; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1012; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1013; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1014; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1015; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1016; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1017; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1018; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1019; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1020; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1021; // @[Mem.scala 73:19:@1120.4]
  wire [31:0] _GEN_1022; // @[Mem.scala 73:19:@1120.4]
  assign _T_1830 = io_mem_addr[31:2]; // @[Mem.scala 65:28:@1111.6]
  assign _T_1834 = _T_1830[7:0]; // @[:@1112.6]
  assign _GEN_0 = 8'h0 == _T_1834 ? io_mem_wdata : memory_0; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_1 = 8'h1 == _T_1834 ? io_mem_wdata : memory_1; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_2 = 8'h2 == _T_1834 ? io_mem_wdata : memory_2; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_3 = 8'h3 == _T_1834 ? io_mem_wdata : memory_3; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_4 = 8'h4 == _T_1834 ? io_mem_wdata : memory_4; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_5 = 8'h5 == _T_1834 ? io_mem_wdata : memory_5; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_6 = 8'h6 == _T_1834 ? io_mem_wdata : memory_6; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_7 = 8'h7 == _T_1834 ? io_mem_wdata : memory_7; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_8 = 8'h8 == _T_1834 ? io_mem_wdata : memory_8; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_9 = 8'h9 == _T_1834 ? io_mem_wdata : memory_9; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_10 = 8'ha == _T_1834 ? io_mem_wdata : memory_10; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_11 = 8'hb == _T_1834 ? io_mem_wdata : memory_11; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_12 = 8'hc == _T_1834 ? io_mem_wdata : memory_12; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_13 = 8'hd == _T_1834 ? io_mem_wdata : memory_13; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_14 = 8'he == _T_1834 ? io_mem_wdata : memory_14; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_15 = 8'hf == _T_1834 ? io_mem_wdata : memory_15; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_16 = 8'h10 == _T_1834 ? io_mem_wdata : memory_16; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_17 = 8'h11 == _T_1834 ? io_mem_wdata : memory_17; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_18 = 8'h12 == _T_1834 ? io_mem_wdata : memory_18; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_19 = 8'h13 == _T_1834 ? io_mem_wdata : memory_19; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_20 = 8'h14 == _T_1834 ? io_mem_wdata : memory_20; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_21 = 8'h15 == _T_1834 ? io_mem_wdata : memory_21; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_22 = 8'h16 == _T_1834 ? io_mem_wdata : memory_22; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_23 = 8'h17 == _T_1834 ? io_mem_wdata : memory_23; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_24 = 8'h18 == _T_1834 ? io_mem_wdata : memory_24; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_25 = 8'h19 == _T_1834 ? io_mem_wdata : memory_25; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_26 = 8'h1a == _T_1834 ? io_mem_wdata : memory_26; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_27 = 8'h1b == _T_1834 ? io_mem_wdata : memory_27; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_28 = 8'h1c == _T_1834 ? io_mem_wdata : memory_28; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_29 = 8'h1d == _T_1834 ? io_mem_wdata : memory_29; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_30 = 8'h1e == _T_1834 ? io_mem_wdata : memory_30; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_31 = 8'h1f == _T_1834 ? io_mem_wdata : memory_31; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_32 = 8'h20 == _T_1834 ? io_mem_wdata : memory_32; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_33 = 8'h21 == _T_1834 ? io_mem_wdata : memory_33; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_34 = 8'h22 == _T_1834 ? io_mem_wdata : memory_34; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_35 = 8'h23 == _T_1834 ? io_mem_wdata : memory_35; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_36 = 8'h24 == _T_1834 ? io_mem_wdata : memory_36; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_37 = 8'h25 == _T_1834 ? io_mem_wdata : memory_37; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_38 = 8'h26 == _T_1834 ? io_mem_wdata : memory_38; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_39 = 8'h27 == _T_1834 ? io_mem_wdata : memory_39; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_40 = 8'h28 == _T_1834 ? io_mem_wdata : memory_40; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_41 = 8'h29 == _T_1834 ? io_mem_wdata : memory_41; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_42 = 8'h2a == _T_1834 ? io_mem_wdata : memory_42; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_43 = 8'h2b == _T_1834 ? io_mem_wdata : memory_43; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_44 = 8'h2c == _T_1834 ? io_mem_wdata : memory_44; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_45 = 8'h2d == _T_1834 ? io_mem_wdata : memory_45; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_46 = 8'h2e == _T_1834 ? io_mem_wdata : memory_46; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_47 = 8'h2f == _T_1834 ? io_mem_wdata : memory_47; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_48 = 8'h30 == _T_1834 ? io_mem_wdata : memory_48; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_49 = 8'h31 == _T_1834 ? io_mem_wdata : memory_49; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_50 = 8'h32 == _T_1834 ? io_mem_wdata : memory_50; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_51 = 8'h33 == _T_1834 ? io_mem_wdata : memory_51; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_52 = 8'h34 == _T_1834 ? io_mem_wdata : memory_52; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_53 = 8'h35 == _T_1834 ? io_mem_wdata : memory_53; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_54 = 8'h36 == _T_1834 ? io_mem_wdata : memory_54; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_55 = 8'h37 == _T_1834 ? io_mem_wdata : memory_55; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_56 = 8'h38 == _T_1834 ? io_mem_wdata : memory_56; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_57 = 8'h39 == _T_1834 ? io_mem_wdata : memory_57; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_58 = 8'h3a == _T_1834 ? io_mem_wdata : memory_58; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_59 = 8'h3b == _T_1834 ? io_mem_wdata : memory_59; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_60 = 8'h3c == _T_1834 ? io_mem_wdata : memory_60; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_61 = 8'h3d == _T_1834 ? io_mem_wdata : memory_61; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_62 = 8'h3e == _T_1834 ? io_mem_wdata : memory_62; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_63 = 8'h3f == _T_1834 ? io_mem_wdata : memory_63; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_64 = 8'h40 == _T_1834 ? io_mem_wdata : memory_64; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_65 = 8'h41 == _T_1834 ? io_mem_wdata : memory_65; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_66 = 8'h42 == _T_1834 ? io_mem_wdata : memory_66; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_67 = 8'h43 == _T_1834 ? io_mem_wdata : memory_67; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_68 = 8'h44 == _T_1834 ? io_mem_wdata : memory_68; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_69 = 8'h45 == _T_1834 ? io_mem_wdata : memory_69; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_70 = 8'h46 == _T_1834 ? io_mem_wdata : memory_70; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_71 = 8'h47 == _T_1834 ? io_mem_wdata : memory_71; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_72 = 8'h48 == _T_1834 ? io_mem_wdata : memory_72; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_73 = 8'h49 == _T_1834 ? io_mem_wdata : memory_73; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_74 = 8'h4a == _T_1834 ? io_mem_wdata : memory_74; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_75 = 8'h4b == _T_1834 ? io_mem_wdata : memory_75; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_76 = 8'h4c == _T_1834 ? io_mem_wdata : memory_76; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_77 = 8'h4d == _T_1834 ? io_mem_wdata : memory_77; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_78 = 8'h4e == _T_1834 ? io_mem_wdata : memory_78; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_79 = 8'h4f == _T_1834 ? io_mem_wdata : memory_79; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_80 = 8'h50 == _T_1834 ? io_mem_wdata : memory_80; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_81 = 8'h51 == _T_1834 ? io_mem_wdata : memory_81; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_82 = 8'h52 == _T_1834 ? io_mem_wdata : memory_82; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_83 = 8'h53 == _T_1834 ? io_mem_wdata : memory_83; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_84 = 8'h54 == _T_1834 ? io_mem_wdata : memory_84; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_85 = 8'h55 == _T_1834 ? io_mem_wdata : memory_85; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_86 = 8'h56 == _T_1834 ? io_mem_wdata : memory_86; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_87 = 8'h57 == _T_1834 ? io_mem_wdata : memory_87; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_88 = 8'h58 == _T_1834 ? io_mem_wdata : memory_88; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_89 = 8'h59 == _T_1834 ? io_mem_wdata : memory_89; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_90 = 8'h5a == _T_1834 ? io_mem_wdata : memory_90; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_91 = 8'h5b == _T_1834 ? io_mem_wdata : memory_91; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_92 = 8'h5c == _T_1834 ? io_mem_wdata : memory_92; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_93 = 8'h5d == _T_1834 ? io_mem_wdata : memory_93; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_94 = 8'h5e == _T_1834 ? io_mem_wdata : memory_94; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_95 = 8'h5f == _T_1834 ? io_mem_wdata : memory_95; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_96 = 8'h60 == _T_1834 ? io_mem_wdata : memory_96; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_97 = 8'h61 == _T_1834 ? io_mem_wdata : memory_97; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_98 = 8'h62 == _T_1834 ? io_mem_wdata : memory_98; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_99 = 8'h63 == _T_1834 ? io_mem_wdata : memory_99; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_100 = 8'h64 == _T_1834 ? io_mem_wdata : memory_100; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_101 = 8'h65 == _T_1834 ? io_mem_wdata : memory_101; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_102 = 8'h66 == _T_1834 ? io_mem_wdata : memory_102; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_103 = 8'h67 == _T_1834 ? io_mem_wdata : memory_103; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_104 = 8'h68 == _T_1834 ? io_mem_wdata : memory_104; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_105 = 8'h69 == _T_1834 ? io_mem_wdata : memory_105; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_106 = 8'h6a == _T_1834 ? io_mem_wdata : memory_106; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_107 = 8'h6b == _T_1834 ? io_mem_wdata : memory_107; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_108 = 8'h6c == _T_1834 ? io_mem_wdata : memory_108; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_109 = 8'h6d == _T_1834 ? io_mem_wdata : memory_109; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_110 = 8'h6e == _T_1834 ? io_mem_wdata : memory_110; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_111 = 8'h6f == _T_1834 ? io_mem_wdata : memory_111; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_112 = 8'h70 == _T_1834 ? io_mem_wdata : memory_112; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_113 = 8'h71 == _T_1834 ? io_mem_wdata : memory_113; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_114 = 8'h72 == _T_1834 ? io_mem_wdata : memory_114; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_115 = 8'h73 == _T_1834 ? io_mem_wdata : memory_115; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_116 = 8'h74 == _T_1834 ? io_mem_wdata : memory_116; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_117 = 8'h75 == _T_1834 ? io_mem_wdata : memory_117; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_118 = 8'h76 == _T_1834 ? io_mem_wdata : memory_118; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_119 = 8'h77 == _T_1834 ? io_mem_wdata : memory_119; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_120 = 8'h78 == _T_1834 ? io_mem_wdata : memory_120; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_121 = 8'h79 == _T_1834 ? io_mem_wdata : memory_121; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_122 = 8'h7a == _T_1834 ? io_mem_wdata : memory_122; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_123 = 8'h7b == _T_1834 ? io_mem_wdata : memory_123; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_124 = 8'h7c == _T_1834 ? io_mem_wdata : memory_124; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_125 = 8'h7d == _T_1834 ? io_mem_wdata : memory_125; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_126 = 8'h7e == _T_1834 ? io_mem_wdata : memory_126; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_127 = 8'h7f == _T_1834 ? io_mem_wdata : memory_127; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_128 = 8'h80 == _T_1834 ? io_mem_wdata : memory_128; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_129 = 8'h81 == _T_1834 ? io_mem_wdata : memory_129; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_130 = 8'h82 == _T_1834 ? io_mem_wdata : memory_130; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_131 = 8'h83 == _T_1834 ? io_mem_wdata : memory_131; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_132 = 8'h84 == _T_1834 ? io_mem_wdata : memory_132; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_133 = 8'h85 == _T_1834 ? io_mem_wdata : memory_133; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_134 = 8'h86 == _T_1834 ? io_mem_wdata : memory_134; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_135 = 8'h87 == _T_1834 ? io_mem_wdata : memory_135; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_136 = 8'h88 == _T_1834 ? io_mem_wdata : memory_136; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_137 = 8'h89 == _T_1834 ? io_mem_wdata : memory_137; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_138 = 8'h8a == _T_1834 ? io_mem_wdata : memory_138; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_139 = 8'h8b == _T_1834 ? io_mem_wdata : memory_139; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_140 = 8'h8c == _T_1834 ? io_mem_wdata : memory_140; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_141 = 8'h8d == _T_1834 ? io_mem_wdata : memory_141; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_142 = 8'h8e == _T_1834 ? io_mem_wdata : memory_142; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_143 = 8'h8f == _T_1834 ? io_mem_wdata : memory_143; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_144 = 8'h90 == _T_1834 ? io_mem_wdata : memory_144; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_145 = 8'h91 == _T_1834 ? io_mem_wdata : memory_145; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_146 = 8'h92 == _T_1834 ? io_mem_wdata : memory_146; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_147 = 8'h93 == _T_1834 ? io_mem_wdata : memory_147; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_148 = 8'h94 == _T_1834 ? io_mem_wdata : memory_148; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_149 = 8'h95 == _T_1834 ? io_mem_wdata : memory_149; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_150 = 8'h96 == _T_1834 ? io_mem_wdata : memory_150; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_151 = 8'h97 == _T_1834 ? io_mem_wdata : memory_151; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_152 = 8'h98 == _T_1834 ? io_mem_wdata : memory_152; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_153 = 8'h99 == _T_1834 ? io_mem_wdata : memory_153; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_154 = 8'h9a == _T_1834 ? io_mem_wdata : memory_154; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_155 = 8'h9b == _T_1834 ? io_mem_wdata : memory_155; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_156 = 8'h9c == _T_1834 ? io_mem_wdata : memory_156; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_157 = 8'h9d == _T_1834 ? io_mem_wdata : memory_157; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_158 = 8'h9e == _T_1834 ? io_mem_wdata : memory_158; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_159 = 8'h9f == _T_1834 ? io_mem_wdata : memory_159; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_160 = 8'ha0 == _T_1834 ? io_mem_wdata : memory_160; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_161 = 8'ha1 == _T_1834 ? io_mem_wdata : memory_161; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_162 = 8'ha2 == _T_1834 ? io_mem_wdata : memory_162; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_163 = 8'ha3 == _T_1834 ? io_mem_wdata : memory_163; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_164 = 8'ha4 == _T_1834 ? io_mem_wdata : memory_164; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_165 = 8'ha5 == _T_1834 ? io_mem_wdata : memory_165; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_166 = 8'ha6 == _T_1834 ? io_mem_wdata : memory_166; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_167 = 8'ha7 == _T_1834 ? io_mem_wdata : memory_167; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_168 = 8'ha8 == _T_1834 ? io_mem_wdata : memory_168; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_169 = 8'ha9 == _T_1834 ? io_mem_wdata : memory_169; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_170 = 8'haa == _T_1834 ? io_mem_wdata : memory_170; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_171 = 8'hab == _T_1834 ? io_mem_wdata : memory_171; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_172 = 8'hac == _T_1834 ? io_mem_wdata : memory_172; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_173 = 8'had == _T_1834 ? io_mem_wdata : memory_173; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_174 = 8'hae == _T_1834 ? io_mem_wdata : memory_174; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_175 = 8'haf == _T_1834 ? io_mem_wdata : memory_175; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_176 = 8'hb0 == _T_1834 ? io_mem_wdata : memory_176; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_177 = 8'hb1 == _T_1834 ? io_mem_wdata : memory_177; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_178 = 8'hb2 == _T_1834 ? io_mem_wdata : memory_178; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_179 = 8'hb3 == _T_1834 ? io_mem_wdata : memory_179; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_180 = 8'hb4 == _T_1834 ? io_mem_wdata : memory_180; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_181 = 8'hb5 == _T_1834 ? io_mem_wdata : memory_181; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_182 = 8'hb6 == _T_1834 ? io_mem_wdata : memory_182; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_183 = 8'hb7 == _T_1834 ? io_mem_wdata : memory_183; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_184 = 8'hb8 == _T_1834 ? io_mem_wdata : memory_184; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_185 = 8'hb9 == _T_1834 ? io_mem_wdata : memory_185; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_186 = 8'hba == _T_1834 ? io_mem_wdata : memory_186; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_187 = 8'hbb == _T_1834 ? io_mem_wdata : memory_187; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_188 = 8'hbc == _T_1834 ? io_mem_wdata : memory_188; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_189 = 8'hbd == _T_1834 ? io_mem_wdata : memory_189; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_190 = 8'hbe == _T_1834 ? io_mem_wdata : memory_190; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_191 = 8'hbf == _T_1834 ? io_mem_wdata : memory_191; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_192 = 8'hc0 == _T_1834 ? io_mem_wdata : memory_192; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_193 = 8'hc1 == _T_1834 ? io_mem_wdata : memory_193; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_194 = 8'hc2 == _T_1834 ? io_mem_wdata : memory_194; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_195 = 8'hc3 == _T_1834 ? io_mem_wdata : memory_195; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_196 = 8'hc4 == _T_1834 ? io_mem_wdata : memory_196; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_197 = 8'hc5 == _T_1834 ? io_mem_wdata : memory_197; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_198 = 8'hc6 == _T_1834 ? io_mem_wdata : memory_198; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_199 = 8'hc7 == _T_1834 ? io_mem_wdata : memory_199; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_200 = 8'hc8 == _T_1834 ? io_mem_wdata : memory_200; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_201 = 8'hc9 == _T_1834 ? io_mem_wdata : memory_201; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_202 = 8'hca == _T_1834 ? io_mem_wdata : memory_202; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_203 = 8'hcb == _T_1834 ? io_mem_wdata : memory_203; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_204 = 8'hcc == _T_1834 ? io_mem_wdata : memory_204; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_205 = 8'hcd == _T_1834 ? io_mem_wdata : memory_205; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_206 = 8'hce == _T_1834 ? io_mem_wdata : memory_206; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_207 = 8'hcf == _T_1834 ? io_mem_wdata : memory_207; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_208 = 8'hd0 == _T_1834 ? io_mem_wdata : memory_208; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_209 = 8'hd1 == _T_1834 ? io_mem_wdata : memory_209; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_210 = 8'hd2 == _T_1834 ? io_mem_wdata : memory_210; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_211 = 8'hd3 == _T_1834 ? io_mem_wdata : memory_211; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_212 = 8'hd4 == _T_1834 ? io_mem_wdata : memory_212; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_213 = 8'hd5 == _T_1834 ? io_mem_wdata : memory_213; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_214 = 8'hd6 == _T_1834 ? io_mem_wdata : memory_214; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_215 = 8'hd7 == _T_1834 ? io_mem_wdata : memory_215; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_216 = 8'hd8 == _T_1834 ? io_mem_wdata : memory_216; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_217 = 8'hd9 == _T_1834 ? io_mem_wdata : memory_217; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_218 = 8'hda == _T_1834 ? io_mem_wdata : memory_218; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_219 = 8'hdb == _T_1834 ? io_mem_wdata : memory_219; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_220 = 8'hdc == _T_1834 ? io_mem_wdata : memory_220; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_221 = 8'hdd == _T_1834 ? io_mem_wdata : memory_221; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_222 = 8'hde == _T_1834 ? io_mem_wdata : memory_222; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_223 = 8'hdf == _T_1834 ? io_mem_wdata : memory_223; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_224 = 8'he0 == _T_1834 ? io_mem_wdata : memory_224; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_225 = 8'he1 == _T_1834 ? io_mem_wdata : memory_225; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_226 = 8'he2 == _T_1834 ? io_mem_wdata : memory_226; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_227 = 8'he3 == _T_1834 ? io_mem_wdata : memory_227; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_228 = 8'he4 == _T_1834 ? io_mem_wdata : memory_228; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_229 = 8'he5 == _T_1834 ? io_mem_wdata : memory_229; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_230 = 8'he6 == _T_1834 ? io_mem_wdata : memory_230; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_231 = 8'he7 == _T_1834 ? io_mem_wdata : memory_231; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_232 = 8'he8 == _T_1834 ? io_mem_wdata : memory_232; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_233 = 8'he9 == _T_1834 ? io_mem_wdata : memory_233; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_234 = 8'hea == _T_1834 ? io_mem_wdata : memory_234; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_235 = 8'heb == _T_1834 ? io_mem_wdata : memory_235; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_236 = 8'hec == _T_1834 ? io_mem_wdata : memory_236; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_237 = 8'hed == _T_1834 ? io_mem_wdata : memory_237; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_238 = 8'hee == _T_1834 ? io_mem_wdata : memory_238; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_239 = 8'hef == _T_1834 ? io_mem_wdata : memory_239; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_240 = 8'hf0 == _T_1834 ? io_mem_wdata : memory_240; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_241 = 8'hf1 == _T_1834 ? io_mem_wdata : memory_241; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_242 = 8'hf2 == _T_1834 ? io_mem_wdata : memory_242; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_243 = 8'hf3 == _T_1834 ? io_mem_wdata : memory_243; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_244 = 8'hf4 == _T_1834 ? io_mem_wdata : memory_244; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_245 = 8'hf5 == _T_1834 ? io_mem_wdata : memory_245; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_246 = 8'hf6 == _T_1834 ? io_mem_wdata : memory_246; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_247 = 8'hf7 == _T_1834 ? io_mem_wdata : memory_247; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_248 = 8'hf8 == _T_1834 ? io_mem_wdata : memory_248; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_249 = 8'hf9 == _T_1834 ? io_mem_wdata : memory_249; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_250 = 8'hfa == _T_1834 ? io_mem_wdata : memory_250; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_251 = 8'hfb == _T_1834 ? io_mem_wdata : memory_251; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_252 = 8'hfc == _T_1834 ? io_mem_wdata : memory_252; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_253 = 8'hfd == _T_1834 ? io_mem_wdata : memory_253; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_254 = 8'hfe == _T_1834 ? io_mem_wdata : memory_254; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_255 = 8'hff == _T_1834 ? io_mem_wdata : memory_255; // @[Mem.scala 65:34:@1113.6]
  assign _GEN_256 = io_mem_wen ? _GEN_0 : memory_0; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_257 = io_mem_wen ? _GEN_1 : memory_1; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_258 = io_mem_wen ? _GEN_2 : memory_2; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_259 = io_mem_wen ? _GEN_3 : memory_3; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_260 = io_mem_wen ? _GEN_4 : memory_4; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_261 = io_mem_wen ? _GEN_5 : memory_5; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_262 = io_mem_wen ? _GEN_6 : memory_6; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_263 = io_mem_wen ? _GEN_7 : memory_7; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_264 = io_mem_wen ? _GEN_8 : memory_8; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_265 = io_mem_wen ? _GEN_9 : memory_9; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_266 = io_mem_wen ? _GEN_10 : memory_10; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_267 = io_mem_wen ? _GEN_11 : memory_11; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_268 = io_mem_wen ? _GEN_12 : memory_12; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_269 = io_mem_wen ? _GEN_13 : memory_13; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_270 = io_mem_wen ? _GEN_14 : memory_14; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_271 = io_mem_wen ? _GEN_15 : memory_15; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_272 = io_mem_wen ? _GEN_16 : memory_16; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_273 = io_mem_wen ? _GEN_17 : memory_17; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_274 = io_mem_wen ? _GEN_18 : memory_18; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_275 = io_mem_wen ? _GEN_19 : memory_19; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_276 = io_mem_wen ? _GEN_20 : memory_20; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_277 = io_mem_wen ? _GEN_21 : memory_21; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_278 = io_mem_wen ? _GEN_22 : memory_22; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_279 = io_mem_wen ? _GEN_23 : memory_23; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_280 = io_mem_wen ? _GEN_24 : memory_24; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_281 = io_mem_wen ? _GEN_25 : memory_25; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_282 = io_mem_wen ? _GEN_26 : memory_26; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_283 = io_mem_wen ? _GEN_27 : memory_27; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_284 = io_mem_wen ? _GEN_28 : memory_28; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_285 = io_mem_wen ? _GEN_29 : memory_29; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_286 = io_mem_wen ? _GEN_30 : memory_30; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_287 = io_mem_wen ? _GEN_31 : memory_31; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_288 = io_mem_wen ? _GEN_32 : memory_32; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_289 = io_mem_wen ? _GEN_33 : memory_33; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_290 = io_mem_wen ? _GEN_34 : memory_34; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_291 = io_mem_wen ? _GEN_35 : memory_35; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_292 = io_mem_wen ? _GEN_36 : memory_36; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_293 = io_mem_wen ? _GEN_37 : memory_37; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_294 = io_mem_wen ? _GEN_38 : memory_38; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_295 = io_mem_wen ? _GEN_39 : memory_39; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_296 = io_mem_wen ? _GEN_40 : memory_40; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_297 = io_mem_wen ? _GEN_41 : memory_41; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_298 = io_mem_wen ? _GEN_42 : memory_42; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_299 = io_mem_wen ? _GEN_43 : memory_43; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_300 = io_mem_wen ? _GEN_44 : memory_44; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_301 = io_mem_wen ? _GEN_45 : memory_45; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_302 = io_mem_wen ? _GEN_46 : memory_46; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_303 = io_mem_wen ? _GEN_47 : memory_47; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_304 = io_mem_wen ? _GEN_48 : memory_48; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_305 = io_mem_wen ? _GEN_49 : memory_49; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_306 = io_mem_wen ? _GEN_50 : memory_50; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_307 = io_mem_wen ? _GEN_51 : memory_51; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_308 = io_mem_wen ? _GEN_52 : memory_52; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_309 = io_mem_wen ? _GEN_53 : memory_53; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_310 = io_mem_wen ? _GEN_54 : memory_54; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_311 = io_mem_wen ? _GEN_55 : memory_55; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_312 = io_mem_wen ? _GEN_56 : memory_56; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_313 = io_mem_wen ? _GEN_57 : memory_57; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_314 = io_mem_wen ? _GEN_58 : memory_58; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_315 = io_mem_wen ? _GEN_59 : memory_59; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_316 = io_mem_wen ? _GEN_60 : memory_60; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_317 = io_mem_wen ? _GEN_61 : memory_61; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_318 = io_mem_wen ? _GEN_62 : memory_62; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_319 = io_mem_wen ? _GEN_63 : memory_63; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_320 = io_mem_wen ? _GEN_64 : memory_64; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_321 = io_mem_wen ? _GEN_65 : memory_65; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_322 = io_mem_wen ? _GEN_66 : memory_66; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_323 = io_mem_wen ? _GEN_67 : memory_67; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_324 = io_mem_wen ? _GEN_68 : memory_68; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_325 = io_mem_wen ? _GEN_69 : memory_69; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_326 = io_mem_wen ? _GEN_70 : memory_70; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_327 = io_mem_wen ? _GEN_71 : memory_71; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_328 = io_mem_wen ? _GEN_72 : memory_72; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_329 = io_mem_wen ? _GEN_73 : memory_73; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_330 = io_mem_wen ? _GEN_74 : memory_74; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_331 = io_mem_wen ? _GEN_75 : memory_75; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_332 = io_mem_wen ? _GEN_76 : memory_76; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_333 = io_mem_wen ? _GEN_77 : memory_77; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_334 = io_mem_wen ? _GEN_78 : memory_78; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_335 = io_mem_wen ? _GEN_79 : memory_79; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_336 = io_mem_wen ? _GEN_80 : memory_80; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_337 = io_mem_wen ? _GEN_81 : memory_81; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_338 = io_mem_wen ? _GEN_82 : memory_82; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_339 = io_mem_wen ? _GEN_83 : memory_83; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_340 = io_mem_wen ? _GEN_84 : memory_84; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_341 = io_mem_wen ? _GEN_85 : memory_85; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_342 = io_mem_wen ? _GEN_86 : memory_86; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_343 = io_mem_wen ? _GEN_87 : memory_87; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_344 = io_mem_wen ? _GEN_88 : memory_88; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_345 = io_mem_wen ? _GEN_89 : memory_89; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_346 = io_mem_wen ? _GEN_90 : memory_90; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_347 = io_mem_wen ? _GEN_91 : memory_91; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_348 = io_mem_wen ? _GEN_92 : memory_92; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_349 = io_mem_wen ? _GEN_93 : memory_93; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_350 = io_mem_wen ? _GEN_94 : memory_94; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_351 = io_mem_wen ? _GEN_95 : memory_95; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_352 = io_mem_wen ? _GEN_96 : memory_96; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_353 = io_mem_wen ? _GEN_97 : memory_97; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_354 = io_mem_wen ? _GEN_98 : memory_98; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_355 = io_mem_wen ? _GEN_99 : memory_99; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_356 = io_mem_wen ? _GEN_100 : memory_100; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_357 = io_mem_wen ? _GEN_101 : memory_101; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_358 = io_mem_wen ? _GEN_102 : memory_102; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_359 = io_mem_wen ? _GEN_103 : memory_103; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_360 = io_mem_wen ? _GEN_104 : memory_104; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_361 = io_mem_wen ? _GEN_105 : memory_105; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_362 = io_mem_wen ? _GEN_106 : memory_106; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_363 = io_mem_wen ? _GEN_107 : memory_107; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_364 = io_mem_wen ? _GEN_108 : memory_108; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_365 = io_mem_wen ? _GEN_109 : memory_109; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_366 = io_mem_wen ? _GEN_110 : memory_110; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_367 = io_mem_wen ? _GEN_111 : memory_111; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_368 = io_mem_wen ? _GEN_112 : memory_112; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_369 = io_mem_wen ? _GEN_113 : memory_113; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_370 = io_mem_wen ? _GEN_114 : memory_114; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_371 = io_mem_wen ? _GEN_115 : memory_115; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_372 = io_mem_wen ? _GEN_116 : memory_116; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_373 = io_mem_wen ? _GEN_117 : memory_117; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_374 = io_mem_wen ? _GEN_118 : memory_118; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_375 = io_mem_wen ? _GEN_119 : memory_119; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_376 = io_mem_wen ? _GEN_120 : memory_120; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_377 = io_mem_wen ? _GEN_121 : memory_121; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_378 = io_mem_wen ? _GEN_122 : memory_122; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_379 = io_mem_wen ? _GEN_123 : memory_123; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_380 = io_mem_wen ? _GEN_124 : memory_124; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_381 = io_mem_wen ? _GEN_125 : memory_125; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_382 = io_mem_wen ? _GEN_126 : memory_126; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_383 = io_mem_wen ? _GEN_127 : memory_127; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_384 = io_mem_wen ? _GEN_128 : memory_128; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_385 = io_mem_wen ? _GEN_129 : memory_129; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_386 = io_mem_wen ? _GEN_130 : memory_130; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_387 = io_mem_wen ? _GEN_131 : memory_131; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_388 = io_mem_wen ? _GEN_132 : memory_132; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_389 = io_mem_wen ? _GEN_133 : memory_133; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_390 = io_mem_wen ? _GEN_134 : memory_134; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_391 = io_mem_wen ? _GEN_135 : memory_135; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_392 = io_mem_wen ? _GEN_136 : memory_136; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_393 = io_mem_wen ? _GEN_137 : memory_137; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_394 = io_mem_wen ? _GEN_138 : memory_138; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_395 = io_mem_wen ? _GEN_139 : memory_139; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_396 = io_mem_wen ? _GEN_140 : memory_140; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_397 = io_mem_wen ? _GEN_141 : memory_141; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_398 = io_mem_wen ? _GEN_142 : memory_142; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_399 = io_mem_wen ? _GEN_143 : memory_143; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_400 = io_mem_wen ? _GEN_144 : memory_144; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_401 = io_mem_wen ? _GEN_145 : memory_145; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_402 = io_mem_wen ? _GEN_146 : memory_146; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_403 = io_mem_wen ? _GEN_147 : memory_147; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_404 = io_mem_wen ? _GEN_148 : memory_148; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_405 = io_mem_wen ? _GEN_149 : memory_149; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_406 = io_mem_wen ? _GEN_150 : memory_150; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_407 = io_mem_wen ? _GEN_151 : memory_151; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_408 = io_mem_wen ? _GEN_152 : memory_152; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_409 = io_mem_wen ? _GEN_153 : memory_153; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_410 = io_mem_wen ? _GEN_154 : memory_154; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_411 = io_mem_wen ? _GEN_155 : memory_155; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_412 = io_mem_wen ? _GEN_156 : memory_156; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_413 = io_mem_wen ? _GEN_157 : memory_157; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_414 = io_mem_wen ? _GEN_158 : memory_158; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_415 = io_mem_wen ? _GEN_159 : memory_159; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_416 = io_mem_wen ? _GEN_160 : memory_160; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_417 = io_mem_wen ? _GEN_161 : memory_161; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_418 = io_mem_wen ? _GEN_162 : memory_162; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_419 = io_mem_wen ? _GEN_163 : memory_163; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_420 = io_mem_wen ? _GEN_164 : memory_164; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_421 = io_mem_wen ? _GEN_165 : memory_165; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_422 = io_mem_wen ? _GEN_166 : memory_166; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_423 = io_mem_wen ? _GEN_167 : memory_167; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_424 = io_mem_wen ? _GEN_168 : memory_168; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_425 = io_mem_wen ? _GEN_169 : memory_169; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_426 = io_mem_wen ? _GEN_170 : memory_170; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_427 = io_mem_wen ? _GEN_171 : memory_171; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_428 = io_mem_wen ? _GEN_172 : memory_172; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_429 = io_mem_wen ? _GEN_173 : memory_173; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_430 = io_mem_wen ? _GEN_174 : memory_174; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_431 = io_mem_wen ? _GEN_175 : memory_175; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_432 = io_mem_wen ? _GEN_176 : memory_176; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_433 = io_mem_wen ? _GEN_177 : memory_177; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_434 = io_mem_wen ? _GEN_178 : memory_178; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_435 = io_mem_wen ? _GEN_179 : memory_179; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_436 = io_mem_wen ? _GEN_180 : memory_180; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_437 = io_mem_wen ? _GEN_181 : memory_181; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_438 = io_mem_wen ? _GEN_182 : memory_182; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_439 = io_mem_wen ? _GEN_183 : memory_183; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_440 = io_mem_wen ? _GEN_184 : memory_184; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_441 = io_mem_wen ? _GEN_185 : memory_185; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_442 = io_mem_wen ? _GEN_186 : memory_186; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_443 = io_mem_wen ? _GEN_187 : memory_187; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_444 = io_mem_wen ? _GEN_188 : memory_188; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_445 = io_mem_wen ? _GEN_189 : memory_189; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_446 = io_mem_wen ? _GEN_190 : memory_190; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_447 = io_mem_wen ? _GEN_191 : memory_191; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_448 = io_mem_wen ? _GEN_192 : memory_192; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_449 = io_mem_wen ? _GEN_193 : memory_193; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_450 = io_mem_wen ? _GEN_194 : memory_194; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_451 = io_mem_wen ? _GEN_195 : memory_195; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_452 = io_mem_wen ? _GEN_196 : memory_196; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_453 = io_mem_wen ? _GEN_197 : memory_197; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_454 = io_mem_wen ? _GEN_198 : memory_198; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_455 = io_mem_wen ? _GEN_199 : memory_199; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_456 = io_mem_wen ? _GEN_200 : memory_200; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_457 = io_mem_wen ? _GEN_201 : memory_201; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_458 = io_mem_wen ? _GEN_202 : memory_202; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_459 = io_mem_wen ? _GEN_203 : memory_203; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_460 = io_mem_wen ? _GEN_204 : memory_204; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_461 = io_mem_wen ? _GEN_205 : memory_205; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_462 = io_mem_wen ? _GEN_206 : memory_206; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_463 = io_mem_wen ? _GEN_207 : memory_207; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_464 = io_mem_wen ? _GEN_208 : memory_208; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_465 = io_mem_wen ? _GEN_209 : memory_209; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_466 = io_mem_wen ? _GEN_210 : memory_210; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_467 = io_mem_wen ? _GEN_211 : memory_211; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_468 = io_mem_wen ? _GEN_212 : memory_212; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_469 = io_mem_wen ? _GEN_213 : memory_213; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_470 = io_mem_wen ? _GEN_214 : memory_214; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_471 = io_mem_wen ? _GEN_215 : memory_215; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_472 = io_mem_wen ? _GEN_216 : memory_216; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_473 = io_mem_wen ? _GEN_217 : memory_217; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_474 = io_mem_wen ? _GEN_218 : memory_218; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_475 = io_mem_wen ? _GEN_219 : memory_219; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_476 = io_mem_wen ? _GEN_220 : memory_220; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_477 = io_mem_wen ? _GEN_221 : memory_221; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_478 = io_mem_wen ? _GEN_222 : memory_222; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_479 = io_mem_wen ? _GEN_223 : memory_223; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_480 = io_mem_wen ? _GEN_224 : memory_224; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_481 = io_mem_wen ? _GEN_225 : memory_225; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_482 = io_mem_wen ? _GEN_226 : memory_226; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_483 = io_mem_wen ? _GEN_227 : memory_227; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_484 = io_mem_wen ? _GEN_228 : memory_228; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_485 = io_mem_wen ? _GEN_229 : memory_229; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_486 = io_mem_wen ? _GEN_230 : memory_230; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_487 = io_mem_wen ? _GEN_231 : memory_231; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_488 = io_mem_wen ? _GEN_232 : memory_232; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_489 = io_mem_wen ? _GEN_233 : memory_233; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_490 = io_mem_wen ? _GEN_234 : memory_234; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_491 = io_mem_wen ? _GEN_235 : memory_235; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_492 = io_mem_wen ? _GEN_236 : memory_236; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_493 = io_mem_wen ? _GEN_237 : memory_237; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_494 = io_mem_wen ? _GEN_238 : memory_238; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_495 = io_mem_wen ? _GEN_239 : memory_239; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_496 = io_mem_wen ? _GEN_240 : memory_240; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_497 = io_mem_wen ? _GEN_241 : memory_241; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_498 = io_mem_wen ? _GEN_242 : memory_242; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_499 = io_mem_wen ? _GEN_243 : memory_243; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_500 = io_mem_wen ? _GEN_244 : memory_244; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_501 = io_mem_wen ? _GEN_245 : memory_245; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_502 = io_mem_wen ? _GEN_246 : memory_246; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_503 = io_mem_wen ? _GEN_247 : memory_247; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_504 = io_mem_wen ? _GEN_248 : memory_248; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_505 = io_mem_wen ? _GEN_249 : memory_249; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_506 = io_mem_wen ? _GEN_250 : memory_250; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_507 = io_mem_wen ? _GEN_251 : memory_251; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_508 = io_mem_wen ? _GEN_252 : memory_252; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_509 = io_mem_wen ? _GEN_253 : memory_253; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_510 = io_mem_wen ? _GEN_254 : memory_254; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_511 = io_mem_wen ? _GEN_255 : memory_255; // @[Mem.scala 64:23:@1110.4]
  assign _GEN_513 = 8'h1 == _T_1834 ? memory_1 : memory_0; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_514 = 8'h2 == _T_1834 ? memory_2 : _GEN_513; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_515 = 8'h3 == _T_1834 ? memory_3 : _GEN_514; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_516 = 8'h4 == _T_1834 ? memory_4 : _GEN_515; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_517 = 8'h5 == _T_1834 ? memory_5 : _GEN_516; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_518 = 8'h6 == _T_1834 ? memory_6 : _GEN_517; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_519 = 8'h7 == _T_1834 ? memory_7 : _GEN_518; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_520 = 8'h8 == _T_1834 ? memory_8 : _GEN_519; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_521 = 8'h9 == _T_1834 ? memory_9 : _GEN_520; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_522 = 8'ha == _T_1834 ? memory_10 : _GEN_521; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_523 = 8'hb == _T_1834 ? memory_11 : _GEN_522; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_524 = 8'hc == _T_1834 ? memory_12 : _GEN_523; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_525 = 8'hd == _T_1834 ? memory_13 : _GEN_524; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_526 = 8'he == _T_1834 ? memory_14 : _GEN_525; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_527 = 8'hf == _T_1834 ? memory_15 : _GEN_526; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_528 = 8'h10 == _T_1834 ? memory_16 : _GEN_527; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_529 = 8'h11 == _T_1834 ? memory_17 : _GEN_528; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_530 = 8'h12 == _T_1834 ? memory_18 : _GEN_529; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_531 = 8'h13 == _T_1834 ? memory_19 : _GEN_530; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_532 = 8'h14 == _T_1834 ? memory_20 : _GEN_531; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_533 = 8'h15 == _T_1834 ? memory_21 : _GEN_532; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_534 = 8'h16 == _T_1834 ? memory_22 : _GEN_533; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_535 = 8'h17 == _T_1834 ? memory_23 : _GEN_534; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_536 = 8'h18 == _T_1834 ? memory_24 : _GEN_535; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_537 = 8'h19 == _T_1834 ? memory_25 : _GEN_536; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_538 = 8'h1a == _T_1834 ? memory_26 : _GEN_537; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_539 = 8'h1b == _T_1834 ? memory_27 : _GEN_538; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_540 = 8'h1c == _T_1834 ? memory_28 : _GEN_539; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_541 = 8'h1d == _T_1834 ? memory_29 : _GEN_540; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_542 = 8'h1e == _T_1834 ? memory_30 : _GEN_541; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_543 = 8'h1f == _T_1834 ? memory_31 : _GEN_542; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_544 = 8'h20 == _T_1834 ? memory_32 : _GEN_543; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_545 = 8'h21 == _T_1834 ? memory_33 : _GEN_544; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_546 = 8'h22 == _T_1834 ? memory_34 : _GEN_545; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_547 = 8'h23 == _T_1834 ? memory_35 : _GEN_546; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_548 = 8'h24 == _T_1834 ? memory_36 : _GEN_547; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_549 = 8'h25 == _T_1834 ? memory_37 : _GEN_548; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_550 = 8'h26 == _T_1834 ? memory_38 : _GEN_549; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_551 = 8'h27 == _T_1834 ? memory_39 : _GEN_550; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_552 = 8'h28 == _T_1834 ? memory_40 : _GEN_551; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_553 = 8'h29 == _T_1834 ? memory_41 : _GEN_552; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_554 = 8'h2a == _T_1834 ? memory_42 : _GEN_553; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_555 = 8'h2b == _T_1834 ? memory_43 : _GEN_554; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_556 = 8'h2c == _T_1834 ? memory_44 : _GEN_555; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_557 = 8'h2d == _T_1834 ? memory_45 : _GEN_556; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_558 = 8'h2e == _T_1834 ? memory_46 : _GEN_557; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_559 = 8'h2f == _T_1834 ? memory_47 : _GEN_558; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_560 = 8'h30 == _T_1834 ? memory_48 : _GEN_559; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_561 = 8'h31 == _T_1834 ? memory_49 : _GEN_560; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_562 = 8'h32 == _T_1834 ? memory_50 : _GEN_561; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_563 = 8'h33 == _T_1834 ? memory_51 : _GEN_562; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_564 = 8'h34 == _T_1834 ? memory_52 : _GEN_563; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_565 = 8'h35 == _T_1834 ? memory_53 : _GEN_564; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_566 = 8'h36 == _T_1834 ? memory_54 : _GEN_565; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_567 = 8'h37 == _T_1834 ? memory_55 : _GEN_566; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_568 = 8'h38 == _T_1834 ? memory_56 : _GEN_567; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_569 = 8'h39 == _T_1834 ? memory_57 : _GEN_568; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_570 = 8'h3a == _T_1834 ? memory_58 : _GEN_569; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_571 = 8'h3b == _T_1834 ? memory_59 : _GEN_570; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_572 = 8'h3c == _T_1834 ? memory_60 : _GEN_571; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_573 = 8'h3d == _T_1834 ? memory_61 : _GEN_572; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_574 = 8'h3e == _T_1834 ? memory_62 : _GEN_573; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_575 = 8'h3f == _T_1834 ? memory_63 : _GEN_574; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_576 = 8'h40 == _T_1834 ? memory_64 : _GEN_575; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_577 = 8'h41 == _T_1834 ? memory_65 : _GEN_576; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_578 = 8'h42 == _T_1834 ? memory_66 : _GEN_577; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_579 = 8'h43 == _T_1834 ? memory_67 : _GEN_578; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_580 = 8'h44 == _T_1834 ? memory_68 : _GEN_579; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_581 = 8'h45 == _T_1834 ? memory_69 : _GEN_580; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_582 = 8'h46 == _T_1834 ? memory_70 : _GEN_581; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_583 = 8'h47 == _T_1834 ? memory_71 : _GEN_582; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_584 = 8'h48 == _T_1834 ? memory_72 : _GEN_583; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_585 = 8'h49 == _T_1834 ? memory_73 : _GEN_584; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_586 = 8'h4a == _T_1834 ? memory_74 : _GEN_585; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_587 = 8'h4b == _T_1834 ? memory_75 : _GEN_586; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_588 = 8'h4c == _T_1834 ? memory_76 : _GEN_587; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_589 = 8'h4d == _T_1834 ? memory_77 : _GEN_588; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_590 = 8'h4e == _T_1834 ? memory_78 : _GEN_589; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_591 = 8'h4f == _T_1834 ? memory_79 : _GEN_590; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_592 = 8'h50 == _T_1834 ? memory_80 : _GEN_591; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_593 = 8'h51 == _T_1834 ? memory_81 : _GEN_592; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_594 = 8'h52 == _T_1834 ? memory_82 : _GEN_593; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_595 = 8'h53 == _T_1834 ? memory_83 : _GEN_594; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_596 = 8'h54 == _T_1834 ? memory_84 : _GEN_595; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_597 = 8'h55 == _T_1834 ? memory_85 : _GEN_596; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_598 = 8'h56 == _T_1834 ? memory_86 : _GEN_597; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_599 = 8'h57 == _T_1834 ? memory_87 : _GEN_598; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_600 = 8'h58 == _T_1834 ? memory_88 : _GEN_599; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_601 = 8'h59 == _T_1834 ? memory_89 : _GEN_600; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_602 = 8'h5a == _T_1834 ? memory_90 : _GEN_601; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_603 = 8'h5b == _T_1834 ? memory_91 : _GEN_602; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_604 = 8'h5c == _T_1834 ? memory_92 : _GEN_603; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_605 = 8'h5d == _T_1834 ? memory_93 : _GEN_604; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_606 = 8'h5e == _T_1834 ? memory_94 : _GEN_605; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_607 = 8'h5f == _T_1834 ? memory_95 : _GEN_606; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_608 = 8'h60 == _T_1834 ? memory_96 : _GEN_607; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_609 = 8'h61 == _T_1834 ? memory_97 : _GEN_608; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_610 = 8'h62 == _T_1834 ? memory_98 : _GEN_609; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_611 = 8'h63 == _T_1834 ? memory_99 : _GEN_610; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_612 = 8'h64 == _T_1834 ? memory_100 : _GEN_611; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_613 = 8'h65 == _T_1834 ? memory_101 : _GEN_612; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_614 = 8'h66 == _T_1834 ? memory_102 : _GEN_613; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_615 = 8'h67 == _T_1834 ? memory_103 : _GEN_614; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_616 = 8'h68 == _T_1834 ? memory_104 : _GEN_615; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_617 = 8'h69 == _T_1834 ? memory_105 : _GEN_616; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_618 = 8'h6a == _T_1834 ? memory_106 : _GEN_617; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_619 = 8'h6b == _T_1834 ? memory_107 : _GEN_618; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_620 = 8'h6c == _T_1834 ? memory_108 : _GEN_619; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_621 = 8'h6d == _T_1834 ? memory_109 : _GEN_620; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_622 = 8'h6e == _T_1834 ? memory_110 : _GEN_621; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_623 = 8'h6f == _T_1834 ? memory_111 : _GEN_622; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_624 = 8'h70 == _T_1834 ? memory_112 : _GEN_623; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_625 = 8'h71 == _T_1834 ? memory_113 : _GEN_624; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_626 = 8'h72 == _T_1834 ? memory_114 : _GEN_625; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_627 = 8'h73 == _T_1834 ? memory_115 : _GEN_626; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_628 = 8'h74 == _T_1834 ? memory_116 : _GEN_627; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_629 = 8'h75 == _T_1834 ? memory_117 : _GEN_628; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_630 = 8'h76 == _T_1834 ? memory_118 : _GEN_629; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_631 = 8'h77 == _T_1834 ? memory_119 : _GEN_630; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_632 = 8'h78 == _T_1834 ? memory_120 : _GEN_631; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_633 = 8'h79 == _T_1834 ? memory_121 : _GEN_632; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_634 = 8'h7a == _T_1834 ? memory_122 : _GEN_633; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_635 = 8'h7b == _T_1834 ? memory_123 : _GEN_634; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_636 = 8'h7c == _T_1834 ? memory_124 : _GEN_635; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_637 = 8'h7d == _T_1834 ? memory_125 : _GEN_636; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_638 = 8'h7e == _T_1834 ? memory_126 : _GEN_637; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_639 = 8'h7f == _T_1834 ? memory_127 : _GEN_638; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_640 = 8'h80 == _T_1834 ? memory_128 : _GEN_639; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_641 = 8'h81 == _T_1834 ? memory_129 : _GEN_640; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_642 = 8'h82 == _T_1834 ? memory_130 : _GEN_641; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_643 = 8'h83 == _T_1834 ? memory_131 : _GEN_642; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_644 = 8'h84 == _T_1834 ? memory_132 : _GEN_643; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_645 = 8'h85 == _T_1834 ? memory_133 : _GEN_644; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_646 = 8'h86 == _T_1834 ? memory_134 : _GEN_645; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_647 = 8'h87 == _T_1834 ? memory_135 : _GEN_646; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_648 = 8'h88 == _T_1834 ? memory_136 : _GEN_647; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_649 = 8'h89 == _T_1834 ? memory_137 : _GEN_648; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_650 = 8'h8a == _T_1834 ? memory_138 : _GEN_649; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_651 = 8'h8b == _T_1834 ? memory_139 : _GEN_650; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_652 = 8'h8c == _T_1834 ? memory_140 : _GEN_651; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_653 = 8'h8d == _T_1834 ? memory_141 : _GEN_652; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_654 = 8'h8e == _T_1834 ? memory_142 : _GEN_653; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_655 = 8'h8f == _T_1834 ? memory_143 : _GEN_654; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_656 = 8'h90 == _T_1834 ? memory_144 : _GEN_655; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_657 = 8'h91 == _T_1834 ? memory_145 : _GEN_656; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_658 = 8'h92 == _T_1834 ? memory_146 : _GEN_657; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_659 = 8'h93 == _T_1834 ? memory_147 : _GEN_658; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_660 = 8'h94 == _T_1834 ? memory_148 : _GEN_659; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_661 = 8'h95 == _T_1834 ? memory_149 : _GEN_660; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_662 = 8'h96 == _T_1834 ? memory_150 : _GEN_661; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_663 = 8'h97 == _T_1834 ? memory_151 : _GEN_662; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_664 = 8'h98 == _T_1834 ? memory_152 : _GEN_663; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_665 = 8'h99 == _T_1834 ? memory_153 : _GEN_664; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_666 = 8'h9a == _T_1834 ? memory_154 : _GEN_665; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_667 = 8'h9b == _T_1834 ? memory_155 : _GEN_666; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_668 = 8'h9c == _T_1834 ? memory_156 : _GEN_667; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_669 = 8'h9d == _T_1834 ? memory_157 : _GEN_668; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_670 = 8'h9e == _T_1834 ? memory_158 : _GEN_669; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_671 = 8'h9f == _T_1834 ? memory_159 : _GEN_670; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_672 = 8'ha0 == _T_1834 ? memory_160 : _GEN_671; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_673 = 8'ha1 == _T_1834 ? memory_161 : _GEN_672; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_674 = 8'ha2 == _T_1834 ? memory_162 : _GEN_673; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_675 = 8'ha3 == _T_1834 ? memory_163 : _GEN_674; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_676 = 8'ha4 == _T_1834 ? memory_164 : _GEN_675; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_677 = 8'ha5 == _T_1834 ? memory_165 : _GEN_676; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_678 = 8'ha6 == _T_1834 ? memory_166 : _GEN_677; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_679 = 8'ha7 == _T_1834 ? memory_167 : _GEN_678; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_680 = 8'ha8 == _T_1834 ? memory_168 : _GEN_679; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_681 = 8'ha9 == _T_1834 ? memory_169 : _GEN_680; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_682 = 8'haa == _T_1834 ? memory_170 : _GEN_681; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_683 = 8'hab == _T_1834 ? memory_171 : _GEN_682; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_684 = 8'hac == _T_1834 ? memory_172 : _GEN_683; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_685 = 8'had == _T_1834 ? memory_173 : _GEN_684; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_686 = 8'hae == _T_1834 ? memory_174 : _GEN_685; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_687 = 8'haf == _T_1834 ? memory_175 : _GEN_686; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_688 = 8'hb0 == _T_1834 ? memory_176 : _GEN_687; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_689 = 8'hb1 == _T_1834 ? memory_177 : _GEN_688; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_690 = 8'hb2 == _T_1834 ? memory_178 : _GEN_689; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_691 = 8'hb3 == _T_1834 ? memory_179 : _GEN_690; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_692 = 8'hb4 == _T_1834 ? memory_180 : _GEN_691; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_693 = 8'hb5 == _T_1834 ? memory_181 : _GEN_692; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_694 = 8'hb6 == _T_1834 ? memory_182 : _GEN_693; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_695 = 8'hb7 == _T_1834 ? memory_183 : _GEN_694; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_696 = 8'hb8 == _T_1834 ? memory_184 : _GEN_695; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_697 = 8'hb9 == _T_1834 ? memory_185 : _GEN_696; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_698 = 8'hba == _T_1834 ? memory_186 : _GEN_697; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_699 = 8'hbb == _T_1834 ? memory_187 : _GEN_698; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_700 = 8'hbc == _T_1834 ? memory_188 : _GEN_699; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_701 = 8'hbd == _T_1834 ? memory_189 : _GEN_700; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_702 = 8'hbe == _T_1834 ? memory_190 : _GEN_701; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_703 = 8'hbf == _T_1834 ? memory_191 : _GEN_702; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_704 = 8'hc0 == _T_1834 ? memory_192 : _GEN_703; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_705 = 8'hc1 == _T_1834 ? memory_193 : _GEN_704; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_706 = 8'hc2 == _T_1834 ? memory_194 : _GEN_705; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_707 = 8'hc3 == _T_1834 ? memory_195 : _GEN_706; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_708 = 8'hc4 == _T_1834 ? memory_196 : _GEN_707; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_709 = 8'hc5 == _T_1834 ? memory_197 : _GEN_708; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_710 = 8'hc6 == _T_1834 ? memory_198 : _GEN_709; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_711 = 8'hc7 == _T_1834 ? memory_199 : _GEN_710; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_712 = 8'hc8 == _T_1834 ? memory_200 : _GEN_711; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_713 = 8'hc9 == _T_1834 ? memory_201 : _GEN_712; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_714 = 8'hca == _T_1834 ? memory_202 : _GEN_713; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_715 = 8'hcb == _T_1834 ? memory_203 : _GEN_714; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_716 = 8'hcc == _T_1834 ? memory_204 : _GEN_715; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_717 = 8'hcd == _T_1834 ? memory_205 : _GEN_716; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_718 = 8'hce == _T_1834 ? memory_206 : _GEN_717; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_719 = 8'hcf == _T_1834 ? memory_207 : _GEN_718; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_720 = 8'hd0 == _T_1834 ? memory_208 : _GEN_719; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_721 = 8'hd1 == _T_1834 ? memory_209 : _GEN_720; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_722 = 8'hd2 == _T_1834 ? memory_210 : _GEN_721; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_723 = 8'hd3 == _T_1834 ? memory_211 : _GEN_722; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_724 = 8'hd4 == _T_1834 ? memory_212 : _GEN_723; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_725 = 8'hd5 == _T_1834 ? memory_213 : _GEN_724; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_726 = 8'hd6 == _T_1834 ? memory_214 : _GEN_725; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_727 = 8'hd7 == _T_1834 ? memory_215 : _GEN_726; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_728 = 8'hd8 == _T_1834 ? memory_216 : _GEN_727; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_729 = 8'hd9 == _T_1834 ? memory_217 : _GEN_728; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_730 = 8'hda == _T_1834 ? memory_218 : _GEN_729; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_731 = 8'hdb == _T_1834 ? memory_219 : _GEN_730; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_732 = 8'hdc == _T_1834 ? memory_220 : _GEN_731; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_733 = 8'hdd == _T_1834 ? memory_221 : _GEN_732; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_734 = 8'hde == _T_1834 ? memory_222 : _GEN_733; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_735 = 8'hdf == _T_1834 ? memory_223 : _GEN_734; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_736 = 8'he0 == _T_1834 ? memory_224 : _GEN_735; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_737 = 8'he1 == _T_1834 ? memory_225 : _GEN_736; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_738 = 8'he2 == _T_1834 ? memory_226 : _GEN_737; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_739 = 8'he3 == _T_1834 ? memory_227 : _GEN_738; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_740 = 8'he4 == _T_1834 ? memory_228 : _GEN_739; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_741 = 8'he5 == _T_1834 ? memory_229 : _GEN_740; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_742 = 8'he6 == _T_1834 ? memory_230 : _GEN_741; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_743 = 8'he7 == _T_1834 ? memory_231 : _GEN_742; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_744 = 8'he8 == _T_1834 ? memory_232 : _GEN_743; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_745 = 8'he9 == _T_1834 ? memory_233 : _GEN_744; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_746 = 8'hea == _T_1834 ? memory_234 : _GEN_745; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_747 = 8'heb == _T_1834 ? memory_235 : _GEN_746; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_748 = 8'hec == _T_1834 ? memory_236 : _GEN_747; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_749 = 8'hed == _T_1834 ? memory_237 : _GEN_748; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_750 = 8'hee == _T_1834 ? memory_238 : _GEN_749; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_751 = 8'hef == _T_1834 ? memory_239 : _GEN_750; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_752 = 8'hf0 == _T_1834 ? memory_240 : _GEN_751; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_753 = 8'hf1 == _T_1834 ? memory_241 : _GEN_752; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_754 = 8'hf2 == _T_1834 ? memory_242 : _GEN_753; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_755 = 8'hf3 == _T_1834 ? memory_243 : _GEN_754; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_756 = 8'hf4 == _T_1834 ? memory_244 : _GEN_755; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_757 = 8'hf5 == _T_1834 ? memory_245 : _GEN_756; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_758 = 8'hf6 == _T_1834 ? memory_246 : _GEN_757; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_759 = 8'hf7 == _T_1834 ? memory_247 : _GEN_758; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_760 = 8'hf8 == _T_1834 ? memory_248 : _GEN_759; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_761 = 8'hf9 == _T_1834 ? memory_249 : _GEN_760; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_762 = 8'hfa == _T_1834 ? memory_250 : _GEN_761; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_763 = 8'hfb == _T_1834 ? memory_251 : _GEN_762; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_764 = 8'hfc == _T_1834 ? memory_252 : _GEN_763; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_765 = 8'hfd == _T_1834 ? memory_253 : _GEN_764; // @[Mem.scala 69:18:@1117.4]
  assign _GEN_766 = 8'hfe == _T_1834 ? memory_254 : _GEN_765; // @[Mem.scala 69:18:@1117.4]
  assign _T_1840 = io_mem_addr2[31:2]; // @[Mem.scala 73:42:@1118.4]
  assign _T_1844 = _T_1840[7:0]; // @[:@1119.4]
  assign _GEN_769 = 8'h1 == _T_1844 ? memory_1 : memory_0; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_770 = 8'h2 == _T_1844 ? memory_2 : _GEN_769; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_771 = 8'h3 == _T_1844 ? memory_3 : _GEN_770; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_772 = 8'h4 == _T_1844 ? memory_4 : _GEN_771; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_773 = 8'h5 == _T_1844 ? memory_5 : _GEN_772; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_774 = 8'h6 == _T_1844 ? memory_6 : _GEN_773; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_775 = 8'h7 == _T_1844 ? memory_7 : _GEN_774; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_776 = 8'h8 == _T_1844 ? memory_8 : _GEN_775; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_777 = 8'h9 == _T_1844 ? memory_9 : _GEN_776; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_778 = 8'ha == _T_1844 ? memory_10 : _GEN_777; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_779 = 8'hb == _T_1844 ? memory_11 : _GEN_778; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_780 = 8'hc == _T_1844 ? memory_12 : _GEN_779; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_781 = 8'hd == _T_1844 ? memory_13 : _GEN_780; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_782 = 8'he == _T_1844 ? memory_14 : _GEN_781; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_783 = 8'hf == _T_1844 ? memory_15 : _GEN_782; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_784 = 8'h10 == _T_1844 ? memory_16 : _GEN_783; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_785 = 8'h11 == _T_1844 ? memory_17 : _GEN_784; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_786 = 8'h12 == _T_1844 ? memory_18 : _GEN_785; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_787 = 8'h13 == _T_1844 ? memory_19 : _GEN_786; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_788 = 8'h14 == _T_1844 ? memory_20 : _GEN_787; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_789 = 8'h15 == _T_1844 ? memory_21 : _GEN_788; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_790 = 8'h16 == _T_1844 ? memory_22 : _GEN_789; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_791 = 8'h17 == _T_1844 ? memory_23 : _GEN_790; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_792 = 8'h18 == _T_1844 ? memory_24 : _GEN_791; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_793 = 8'h19 == _T_1844 ? memory_25 : _GEN_792; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_794 = 8'h1a == _T_1844 ? memory_26 : _GEN_793; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_795 = 8'h1b == _T_1844 ? memory_27 : _GEN_794; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_796 = 8'h1c == _T_1844 ? memory_28 : _GEN_795; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_797 = 8'h1d == _T_1844 ? memory_29 : _GEN_796; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_798 = 8'h1e == _T_1844 ? memory_30 : _GEN_797; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_799 = 8'h1f == _T_1844 ? memory_31 : _GEN_798; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_800 = 8'h20 == _T_1844 ? memory_32 : _GEN_799; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_801 = 8'h21 == _T_1844 ? memory_33 : _GEN_800; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_802 = 8'h22 == _T_1844 ? memory_34 : _GEN_801; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_803 = 8'h23 == _T_1844 ? memory_35 : _GEN_802; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_804 = 8'h24 == _T_1844 ? memory_36 : _GEN_803; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_805 = 8'h25 == _T_1844 ? memory_37 : _GEN_804; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_806 = 8'h26 == _T_1844 ? memory_38 : _GEN_805; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_807 = 8'h27 == _T_1844 ? memory_39 : _GEN_806; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_808 = 8'h28 == _T_1844 ? memory_40 : _GEN_807; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_809 = 8'h29 == _T_1844 ? memory_41 : _GEN_808; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_810 = 8'h2a == _T_1844 ? memory_42 : _GEN_809; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_811 = 8'h2b == _T_1844 ? memory_43 : _GEN_810; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_812 = 8'h2c == _T_1844 ? memory_44 : _GEN_811; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_813 = 8'h2d == _T_1844 ? memory_45 : _GEN_812; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_814 = 8'h2e == _T_1844 ? memory_46 : _GEN_813; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_815 = 8'h2f == _T_1844 ? memory_47 : _GEN_814; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_816 = 8'h30 == _T_1844 ? memory_48 : _GEN_815; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_817 = 8'h31 == _T_1844 ? memory_49 : _GEN_816; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_818 = 8'h32 == _T_1844 ? memory_50 : _GEN_817; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_819 = 8'h33 == _T_1844 ? memory_51 : _GEN_818; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_820 = 8'h34 == _T_1844 ? memory_52 : _GEN_819; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_821 = 8'h35 == _T_1844 ? memory_53 : _GEN_820; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_822 = 8'h36 == _T_1844 ? memory_54 : _GEN_821; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_823 = 8'h37 == _T_1844 ? memory_55 : _GEN_822; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_824 = 8'h38 == _T_1844 ? memory_56 : _GEN_823; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_825 = 8'h39 == _T_1844 ? memory_57 : _GEN_824; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_826 = 8'h3a == _T_1844 ? memory_58 : _GEN_825; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_827 = 8'h3b == _T_1844 ? memory_59 : _GEN_826; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_828 = 8'h3c == _T_1844 ? memory_60 : _GEN_827; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_829 = 8'h3d == _T_1844 ? memory_61 : _GEN_828; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_830 = 8'h3e == _T_1844 ? memory_62 : _GEN_829; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_831 = 8'h3f == _T_1844 ? memory_63 : _GEN_830; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_832 = 8'h40 == _T_1844 ? memory_64 : _GEN_831; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_833 = 8'h41 == _T_1844 ? memory_65 : _GEN_832; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_834 = 8'h42 == _T_1844 ? memory_66 : _GEN_833; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_835 = 8'h43 == _T_1844 ? memory_67 : _GEN_834; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_836 = 8'h44 == _T_1844 ? memory_68 : _GEN_835; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_837 = 8'h45 == _T_1844 ? memory_69 : _GEN_836; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_838 = 8'h46 == _T_1844 ? memory_70 : _GEN_837; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_839 = 8'h47 == _T_1844 ? memory_71 : _GEN_838; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_840 = 8'h48 == _T_1844 ? memory_72 : _GEN_839; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_841 = 8'h49 == _T_1844 ? memory_73 : _GEN_840; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_842 = 8'h4a == _T_1844 ? memory_74 : _GEN_841; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_843 = 8'h4b == _T_1844 ? memory_75 : _GEN_842; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_844 = 8'h4c == _T_1844 ? memory_76 : _GEN_843; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_845 = 8'h4d == _T_1844 ? memory_77 : _GEN_844; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_846 = 8'h4e == _T_1844 ? memory_78 : _GEN_845; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_847 = 8'h4f == _T_1844 ? memory_79 : _GEN_846; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_848 = 8'h50 == _T_1844 ? memory_80 : _GEN_847; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_849 = 8'h51 == _T_1844 ? memory_81 : _GEN_848; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_850 = 8'h52 == _T_1844 ? memory_82 : _GEN_849; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_851 = 8'h53 == _T_1844 ? memory_83 : _GEN_850; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_852 = 8'h54 == _T_1844 ? memory_84 : _GEN_851; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_853 = 8'h55 == _T_1844 ? memory_85 : _GEN_852; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_854 = 8'h56 == _T_1844 ? memory_86 : _GEN_853; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_855 = 8'h57 == _T_1844 ? memory_87 : _GEN_854; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_856 = 8'h58 == _T_1844 ? memory_88 : _GEN_855; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_857 = 8'h59 == _T_1844 ? memory_89 : _GEN_856; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_858 = 8'h5a == _T_1844 ? memory_90 : _GEN_857; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_859 = 8'h5b == _T_1844 ? memory_91 : _GEN_858; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_860 = 8'h5c == _T_1844 ? memory_92 : _GEN_859; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_861 = 8'h5d == _T_1844 ? memory_93 : _GEN_860; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_862 = 8'h5e == _T_1844 ? memory_94 : _GEN_861; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_863 = 8'h5f == _T_1844 ? memory_95 : _GEN_862; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_864 = 8'h60 == _T_1844 ? memory_96 : _GEN_863; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_865 = 8'h61 == _T_1844 ? memory_97 : _GEN_864; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_866 = 8'h62 == _T_1844 ? memory_98 : _GEN_865; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_867 = 8'h63 == _T_1844 ? memory_99 : _GEN_866; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_868 = 8'h64 == _T_1844 ? memory_100 : _GEN_867; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_869 = 8'h65 == _T_1844 ? memory_101 : _GEN_868; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_870 = 8'h66 == _T_1844 ? memory_102 : _GEN_869; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_871 = 8'h67 == _T_1844 ? memory_103 : _GEN_870; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_872 = 8'h68 == _T_1844 ? memory_104 : _GEN_871; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_873 = 8'h69 == _T_1844 ? memory_105 : _GEN_872; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_874 = 8'h6a == _T_1844 ? memory_106 : _GEN_873; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_875 = 8'h6b == _T_1844 ? memory_107 : _GEN_874; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_876 = 8'h6c == _T_1844 ? memory_108 : _GEN_875; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_877 = 8'h6d == _T_1844 ? memory_109 : _GEN_876; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_878 = 8'h6e == _T_1844 ? memory_110 : _GEN_877; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_879 = 8'h6f == _T_1844 ? memory_111 : _GEN_878; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_880 = 8'h70 == _T_1844 ? memory_112 : _GEN_879; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_881 = 8'h71 == _T_1844 ? memory_113 : _GEN_880; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_882 = 8'h72 == _T_1844 ? memory_114 : _GEN_881; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_883 = 8'h73 == _T_1844 ? memory_115 : _GEN_882; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_884 = 8'h74 == _T_1844 ? memory_116 : _GEN_883; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_885 = 8'h75 == _T_1844 ? memory_117 : _GEN_884; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_886 = 8'h76 == _T_1844 ? memory_118 : _GEN_885; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_887 = 8'h77 == _T_1844 ? memory_119 : _GEN_886; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_888 = 8'h78 == _T_1844 ? memory_120 : _GEN_887; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_889 = 8'h79 == _T_1844 ? memory_121 : _GEN_888; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_890 = 8'h7a == _T_1844 ? memory_122 : _GEN_889; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_891 = 8'h7b == _T_1844 ? memory_123 : _GEN_890; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_892 = 8'h7c == _T_1844 ? memory_124 : _GEN_891; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_893 = 8'h7d == _T_1844 ? memory_125 : _GEN_892; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_894 = 8'h7e == _T_1844 ? memory_126 : _GEN_893; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_895 = 8'h7f == _T_1844 ? memory_127 : _GEN_894; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_896 = 8'h80 == _T_1844 ? memory_128 : _GEN_895; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_897 = 8'h81 == _T_1844 ? memory_129 : _GEN_896; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_898 = 8'h82 == _T_1844 ? memory_130 : _GEN_897; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_899 = 8'h83 == _T_1844 ? memory_131 : _GEN_898; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_900 = 8'h84 == _T_1844 ? memory_132 : _GEN_899; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_901 = 8'h85 == _T_1844 ? memory_133 : _GEN_900; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_902 = 8'h86 == _T_1844 ? memory_134 : _GEN_901; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_903 = 8'h87 == _T_1844 ? memory_135 : _GEN_902; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_904 = 8'h88 == _T_1844 ? memory_136 : _GEN_903; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_905 = 8'h89 == _T_1844 ? memory_137 : _GEN_904; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_906 = 8'h8a == _T_1844 ? memory_138 : _GEN_905; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_907 = 8'h8b == _T_1844 ? memory_139 : _GEN_906; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_908 = 8'h8c == _T_1844 ? memory_140 : _GEN_907; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_909 = 8'h8d == _T_1844 ? memory_141 : _GEN_908; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_910 = 8'h8e == _T_1844 ? memory_142 : _GEN_909; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_911 = 8'h8f == _T_1844 ? memory_143 : _GEN_910; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_912 = 8'h90 == _T_1844 ? memory_144 : _GEN_911; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_913 = 8'h91 == _T_1844 ? memory_145 : _GEN_912; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_914 = 8'h92 == _T_1844 ? memory_146 : _GEN_913; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_915 = 8'h93 == _T_1844 ? memory_147 : _GEN_914; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_916 = 8'h94 == _T_1844 ? memory_148 : _GEN_915; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_917 = 8'h95 == _T_1844 ? memory_149 : _GEN_916; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_918 = 8'h96 == _T_1844 ? memory_150 : _GEN_917; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_919 = 8'h97 == _T_1844 ? memory_151 : _GEN_918; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_920 = 8'h98 == _T_1844 ? memory_152 : _GEN_919; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_921 = 8'h99 == _T_1844 ? memory_153 : _GEN_920; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_922 = 8'h9a == _T_1844 ? memory_154 : _GEN_921; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_923 = 8'h9b == _T_1844 ? memory_155 : _GEN_922; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_924 = 8'h9c == _T_1844 ? memory_156 : _GEN_923; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_925 = 8'h9d == _T_1844 ? memory_157 : _GEN_924; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_926 = 8'h9e == _T_1844 ? memory_158 : _GEN_925; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_927 = 8'h9f == _T_1844 ? memory_159 : _GEN_926; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_928 = 8'ha0 == _T_1844 ? memory_160 : _GEN_927; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_929 = 8'ha1 == _T_1844 ? memory_161 : _GEN_928; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_930 = 8'ha2 == _T_1844 ? memory_162 : _GEN_929; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_931 = 8'ha3 == _T_1844 ? memory_163 : _GEN_930; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_932 = 8'ha4 == _T_1844 ? memory_164 : _GEN_931; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_933 = 8'ha5 == _T_1844 ? memory_165 : _GEN_932; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_934 = 8'ha6 == _T_1844 ? memory_166 : _GEN_933; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_935 = 8'ha7 == _T_1844 ? memory_167 : _GEN_934; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_936 = 8'ha8 == _T_1844 ? memory_168 : _GEN_935; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_937 = 8'ha9 == _T_1844 ? memory_169 : _GEN_936; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_938 = 8'haa == _T_1844 ? memory_170 : _GEN_937; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_939 = 8'hab == _T_1844 ? memory_171 : _GEN_938; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_940 = 8'hac == _T_1844 ? memory_172 : _GEN_939; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_941 = 8'had == _T_1844 ? memory_173 : _GEN_940; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_942 = 8'hae == _T_1844 ? memory_174 : _GEN_941; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_943 = 8'haf == _T_1844 ? memory_175 : _GEN_942; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_944 = 8'hb0 == _T_1844 ? memory_176 : _GEN_943; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_945 = 8'hb1 == _T_1844 ? memory_177 : _GEN_944; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_946 = 8'hb2 == _T_1844 ? memory_178 : _GEN_945; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_947 = 8'hb3 == _T_1844 ? memory_179 : _GEN_946; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_948 = 8'hb4 == _T_1844 ? memory_180 : _GEN_947; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_949 = 8'hb5 == _T_1844 ? memory_181 : _GEN_948; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_950 = 8'hb6 == _T_1844 ? memory_182 : _GEN_949; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_951 = 8'hb7 == _T_1844 ? memory_183 : _GEN_950; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_952 = 8'hb8 == _T_1844 ? memory_184 : _GEN_951; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_953 = 8'hb9 == _T_1844 ? memory_185 : _GEN_952; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_954 = 8'hba == _T_1844 ? memory_186 : _GEN_953; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_955 = 8'hbb == _T_1844 ? memory_187 : _GEN_954; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_956 = 8'hbc == _T_1844 ? memory_188 : _GEN_955; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_957 = 8'hbd == _T_1844 ? memory_189 : _GEN_956; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_958 = 8'hbe == _T_1844 ? memory_190 : _GEN_957; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_959 = 8'hbf == _T_1844 ? memory_191 : _GEN_958; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_960 = 8'hc0 == _T_1844 ? memory_192 : _GEN_959; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_961 = 8'hc1 == _T_1844 ? memory_193 : _GEN_960; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_962 = 8'hc2 == _T_1844 ? memory_194 : _GEN_961; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_963 = 8'hc3 == _T_1844 ? memory_195 : _GEN_962; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_964 = 8'hc4 == _T_1844 ? memory_196 : _GEN_963; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_965 = 8'hc5 == _T_1844 ? memory_197 : _GEN_964; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_966 = 8'hc6 == _T_1844 ? memory_198 : _GEN_965; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_967 = 8'hc7 == _T_1844 ? memory_199 : _GEN_966; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_968 = 8'hc8 == _T_1844 ? memory_200 : _GEN_967; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_969 = 8'hc9 == _T_1844 ? memory_201 : _GEN_968; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_970 = 8'hca == _T_1844 ? memory_202 : _GEN_969; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_971 = 8'hcb == _T_1844 ? memory_203 : _GEN_970; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_972 = 8'hcc == _T_1844 ? memory_204 : _GEN_971; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_973 = 8'hcd == _T_1844 ? memory_205 : _GEN_972; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_974 = 8'hce == _T_1844 ? memory_206 : _GEN_973; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_975 = 8'hcf == _T_1844 ? memory_207 : _GEN_974; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_976 = 8'hd0 == _T_1844 ? memory_208 : _GEN_975; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_977 = 8'hd1 == _T_1844 ? memory_209 : _GEN_976; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_978 = 8'hd2 == _T_1844 ? memory_210 : _GEN_977; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_979 = 8'hd3 == _T_1844 ? memory_211 : _GEN_978; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_980 = 8'hd4 == _T_1844 ? memory_212 : _GEN_979; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_981 = 8'hd5 == _T_1844 ? memory_213 : _GEN_980; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_982 = 8'hd6 == _T_1844 ? memory_214 : _GEN_981; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_983 = 8'hd7 == _T_1844 ? memory_215 : _GEN_982; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_984 = 8'hd8 == _T_1844 ? memory_216 : _GEN_983; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_985 = 8'hd9 == _T_1844 ? memory_217 : _GEN_984; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_986 = 8'hda == _T_1844 ? memory_218 : _GEN_985; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_987 = 8'hdb == _T_1844 ? memory_219 : _GEN_986; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_988 = 8'hdc == _T_1844 ? memory_220 : _GEN_987; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_989 = 8'hdd == _T_1844 ? memory_221 : _GEN_988; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_990 = 8'hde == _T_1844 ? memory_222 : _GEN_989; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_991 = 8'hdf == _T_1844 ? memory_223 : _GEN_990; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_992 = 8'he0 == _T_1844 ? memory_224 : _GEN_991; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_993 = 8'he1 == _T_1844 ? memory_225 : _GEN_992; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_994 = 8'he2 == _T_1844 ? memory_226 : _GEN_993; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_995 = 8'he3 == _T_1844 ? memory_227 : _GEN_994; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_996 = 8'he4 == _T_1844 ? memory_228 : _GEN_995; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_997 = 8'he5 == _T_1844 ? memory_229 : _GEN_996; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_998 = 8'he6 == _T_1844 ? memory_230 : _GEN_997; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_999 = 8'he7 == _T_1844 ? memory_231 : _GEN_998; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1000 = 8'he8 == _T_1844 ? memory_232 : _GEN_999; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1001 = 8'he9 == _T_1844 ? memory_233 : _GEN_1000; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1002 = 8'hea == _T_1844 ? memory_234 : _GEN_1001; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1003 = 8'heb == _T_1844 ? memory_235 : _GEN_1002; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1004 = 8'hec == _T_1844 ? memory_236 : _GEN_1003; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1005 = 8'hed == _T_1844 ? memory_237 : _GEN_1004; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1006 = 8'hee == _T_1844 ? memory_238 : _GEN_1005; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1007 = 8'hef == _T_1844 ? memory_239 : _GEN_1006; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1008 = 8'hf0 == _T_1844 ? memory_240 : _GEN_1007; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1009 = 8'hf1 == _T_1844 ? memory_241 : _GEN_1008; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1010 = 8'hf2 == _T_1844 ? memory_242 : _GEN_1009; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1011 = 8'hf3 == _T_1844 ? memory_243 : _GEN_1010; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1012 = 8'hf4 == _T_1844 ? memory_244 : _GEN_1011; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1013 = 8'hf5 == _T_1844 ? memory_245 : _GEN_1012; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1014 = 8'hf6 == _T_1844 ? memory_246 : _GEN_1013; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1015 = 8'hf7 == _T_1844 ? memory_247 : _GEN_1014; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1016 = 8'hf8 == _T_1844 ? memory_248 : _GEN_1015; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1017 = 8'hf9 == _T_1844 ? memory_249 : _GEN_1016; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1018 = 8'hfa == _T_1844 ? memory_250 : _GEN_1017; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1019 = 8'hfb == _T_1844 ? memory_251 : _GEN_1018; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1020 = 8'hfc == _T_1844 ? memory_252 : _GEN_1019; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1021 = 8'hfd == _T_1844 ? memory_253 : _GEN_1020; // @[Mem.scala 73:19:@1120.4]
  assign _GEN_1022 = 8'hfe == _T_1844 ? memory_254 : _GEN_1021; // @[Mem.scala 73:19:@1120.4]
  assign io_mem_rdata = 8'hff == _T_1834 ? memory_255 : _GEN_766; // @[Mem.scala 69:18:@1117.4]
  assign io_mem_rdata2 = 8'hff == _T_1844 ? memory_255 : _GEN_1022; // @[Mem.scala 73:19:@1120.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  memory_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  memory_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  memory_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  memory_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  memory_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  memory_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  memory_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  memory_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  memory_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  memory_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  memory_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  memory_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  memory_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  memory_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  memory_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  memory_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  memory_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  memory_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  memory_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  memory_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  memory_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  memory_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  memory_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  memory_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  memory_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  memory_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  memory_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  memory_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  memory_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  memory_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  memory_30 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  memory_31 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  memory_32 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  memory_33 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  memory_34 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  memory_35 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  memory_36 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  memory_37 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  memory_38 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  memory_39 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  memory_40 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  memory_41 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  memory_42 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  memory_43 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  memory_44 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  memory_45 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  memory_46 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  memory_47 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  memory_48 = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  memory_49 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  memory_50 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  memory_51 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  memory_52 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  memory_53 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  memory_54 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  memory_55 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  memory_56 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  memory_57 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  memory_58 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  memory_59 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  memory_60 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  memory_61 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  memory_62 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  memory_63 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  memory_64 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  memory_65 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  memory_66 = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  memory_67 = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  memory_68 = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  memory_69 = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  memory_70 = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  memory_71 = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  memory_72 = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  memory_73 = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  memory_74 = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  memory_75 = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  memory_76 = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  memory_77 = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  memory_78 = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  memory_79 = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  memory_80 = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  memory_81 = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  memory_82 = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  memory_83 = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  memory_84 = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  memory_85 = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  memory_86 = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  memory_87 = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  memory_88 = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  memory_89 = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  memory_90 = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  memory_91 = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  memory_92 = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  memory_93 = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  memory_94 = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  memory_95 = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  memory_96 = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  memory_97 = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  memory_98 = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  memory_99 = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  memory_100 = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  memory_101 = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  memory_102 = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  memory_103 = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  memory_104 = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  memory_105 = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  memory_106 = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  memory_107 = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  memory_108 = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  memory_109 = _RAND_109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  memory_110 = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  memory_111 = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  memory_112 = _RAND_112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  memory_113 = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  memory_114 = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  memory_115 = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  memory_116 = _RAND_116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  memory_117 = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  memory_118 = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  memory_119 = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  memory_120 = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  memory_121 = _RAND_121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  memory_122 = _RAND_122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  memory_123 = _RAND_123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  memory_124 = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  memory_125 = _RAND_125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  memory_126 = _RAND_126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  memory_127 = _RAND_127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  memory_128 = _RAND_128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  memory_129 = _RAND_129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  memory_130 = _RAND_130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  memory_131 = _RAND_131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  memory_132 = _RAND_132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  memory_133 = _RAND_133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  memory_134 = _RAND_134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  memory_135 = _RAND_135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  memory_136 = _RAND_136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  memory_137 = _RAND_137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  memory_138 = _RAND_138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  memory_139 = _RAND_139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  memory_140 = _RAND_140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  memory_141 = _RAND_141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  memory_142 = _RAND_142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  memory_143 = _RAND_143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  memory_144 = _RAND_144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  memory_145 = _RAND_145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  memory_146 = _RAND_146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  memory_147 = _RAND_147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  memory_148 = _RAND_148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  memory_149 = _RAND_149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  memory_150 = _RAND_150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  memory_151 = _RAND_151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  memory_152 = _RAND_152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  memory_153 = _RAND_153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  memory_154 = _RAND_154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  memory_155 = _RAND_155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  memory_156 = _RAND_156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  memory_157 = _RAND_157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  memory_158 = _RAND_158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  memory_159 = _RAND_159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  memory_160 = _RAND_160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  memory_161 = _RAND_161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  memory_162 = _RAND_162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  memory_163 = _RAND_163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  memory_164 = _RAND_164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  memory_165 = _RAND_165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  memory_166 = _RAND_166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  memory_167 = _RAND_167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  memory_168 = _RAND_168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  memory_169 = _RAND_169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  memory_170 = _RAND_170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  memory_171 = _RAND_171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  memory_172 = _RAND_172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  memory_173 = _RAND_173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  memory_174 = _RAND_174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  memory_175 = _RAND_175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  memory_176 = _RAND_176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  memory_177 = _RAND_177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  memory_178 = _RAND_178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  memory_179 = _RAND_179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  memory_180 = _RAND_180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  memory_181 = _RAND_181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  memory_182 = _RAND_182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  memory_183 = _RAND_183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  memory_184 = _RAND_184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  memory_185 = _RAND_185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  memory_186 = _RAND_186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  memory_187 = _RAND_187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  memory_188 = _RAND_188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  memory_189 = _RAND_189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  memory_190 = _RAND_190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  memory_191 = _RAND_191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  memory_192 = _RAND_192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  memory_193 = _RAND_193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  memory_194 = _RAND_194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  memory_195 = _RAND_195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  memory_196 = _RAND_196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  memory_197 = _RAND_197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  memory_198 = _RAND_198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  memory_199 = _RAND_199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  memory_200 = _RAND_200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  memory_201 = _RAND_201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  memory_202 = _RAND_202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  memory_203 = _RAND_203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  memory_204 = _RAND_204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  memory_205 = _RAND_205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  memory_206 = _RAND_206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  memory_207 = _RAND_207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  memory_208 = _RAND_208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  memory_209 = _RAND_209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  memory_210 = _RAND_210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  memory_211 = _RAND_211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  memory_212 = _RAND_212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  memory_213 = _RAND_213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  memory_214 = _RAND_214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  memory_215 = _RAND_215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  memory_216 = _RAND_216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  memory_217 = _RAND_217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  memory_218 = _RAND_218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  memory_219 = _RAND_219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  memory_220 = _RAND_220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  memory_221 = _RAND_221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  memory_222 = _RAND_222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  memory_223 = _RAND_223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  memory_224 = _RAND_224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  memory_225 = _RAND_225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  memory_226 = _RAND_226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  memory_227 = _RAND_227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  memory_228 = _RAND_228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  memory_229 = _RAND_229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  memory_230 = _RAND_230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  memory_231 = _RAND_231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  memory_232 = _RAND_232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  memory_233 = _RAND_233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  memory_234 = _RAND_234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  memory_235 = _RAND_235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  memory_236 = _RAND_236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  memory_237 = _RAND_237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  memory_238 = _RAND_238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  memory_239 = _RAND_239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  memory_240 = _RAND_240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  memory_241 = _RAND_241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  memory_242 = _RAND_242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  memory_243 = _RAND_243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  memory_244 = _RAND_244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  memory_245 = _RAND_245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  memory_246 = _RAND_246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  memory_247 = _RAND_247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  memory_248 = _RAND_248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  memory_249 = _RAND_249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  memory_250 = _RAND_250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  memory_251 = _RAND_251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  memory_252 = _RAND_252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  memory_253 = _RAND_253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  memory_254 = _RAND_254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  memory_255 = _RAND_255[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      memory_0 <= 32'h201d03fc;
    end else begin
      if (io_mem_wen) begin
        if (8'h0 == _T_1834) begin
          memory_0 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_1 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h1 == _T_1834) begin
          memory_1 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_2 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h2 == _T_1834) begin
          memory_2 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_3 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h3 == _T_1834) begin
          memory_3 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_4 <= 32'h27bdffd8;
    end else begin
      if (io_mem_wen) begin
        if (8'h4 == _T_1834) begin
          memory_4 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_5 <= 32'hafbf0024;
    end else begin
      if (io_mem_wen) begin
        if (8'h5 == _T_1834) begin
          memory_5 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_6 <= 32'hafbe0020;
    end else begin
      if (io_mem_wen) begin
        if (8'h6 == _T_1834) begin
          memory_6 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_7 <= 32'h3a0f025;
    end else begin
      if (io_mem_wen) begin
        if (8'h7 == _T_1834) begin
          memory_7 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_8 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h8 == _T_1834) begin
          memory_8 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_9 <= 32'hac400350;
    end else begin
      if (io_mem_wen) begin
        if (8'h9 == _T_1834) begin
          memory_9 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_10 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'ha == _T_1834) begin
          memory_10 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_11 <= 32'hac400354;
    end else begin
      if (io_mem_wen) begin
        if (8'hb == _T_1834) begin
          memory_11 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_12 <= 32'h24040f3e;
    end else begin
      if (io_mem_wen) begin
        if (8'hc == _T_1834) begin
          memory_12 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_13 <= 32'hc000076;
    end else begin
      if (io_mem_wen) begin
        if (8'hd == _T_1834) begin
          memory_13 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_14 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'he == _T_1834) begin
          memory_14 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_15 <= 32'hc0000af;
    end else begin
      if (io_mem_wen) begin
        if (8'hf == _T_1834) begin
          memory_15 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_16 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h10 == _T_1834) begin
          memory_16 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_17 <= 32'hafc2001c;
    end else begin
      if (io_mem_wen) begin
        if (8'h11 == _T_1834) begin
          memory_17 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_18 <= 32'h8fc3001c;
    end else begin
      if (io_mem_wen) begin
        if (8'h12 == _T_1834) begin
          memory_18 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_19 <= 32'h2402000a;
    end else begin
      if (io_mem_wen) begin
        if (8'h13 == _T_1834) begin
          memory_19 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_20 <= 32'h10620005;
    end else begin
      if (io_mem_wen) begin
        if (8'h14 == _T_1834) begin
          memory_20 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_21 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h15 == _T_1834) begin
          memory_21 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_22 <= 32'h8fc3001c;
    end else begin
      if (io_mem_wen) begin
        if (8'h16 == _T_1834) begin
          memory_22 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_23 <= 32'h2402000d;
    end else begin
      if (io_mem_wen) begin
        if (8'h17 == _T_1834) begin
          memory_23 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_24 <= 32'h1462000b;
    end else begin
      if (io_mem_wen) begin
        if (8'h18 == _T_1834) begin
          memory_24 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_25 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h19 == _T_1834) begin
          memory_25 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_26 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h1a == _T_1834) begin
          memory_26 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_27 <= 32'hac400350;
    end else begin
      if (io_mem_wen) begin
        if (8'h1b == _T_1834) begin
          memory_27 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_28 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h1c == _T_1834) begin
          memory_28 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_29 <= 32'h8c420354;
    end else begin
      if (io_mem_wen) begin
        if (8'h1d == _T_1834) begin
          memory_29 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_30 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h1e == _T_1834) begin
          memory_30 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_31 <= 32'h24430001;
    end else begin
      if (io_mem_wen) begin
        if (8'h1f == _T_1834) begin
          memory_31 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_32 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h20 == _T_1834) begin
          memory_32 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_33 <= 32'hac430354;
    end else begin
      if (io_mem_wen) begin
        if (8'h21 == _T_1834) begin
          memory_33 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_34 <= 32'h10000051;
    end else begin
      if (io_mem_wen) begin
        if (8'h22 == _T_1834) begin
          memory_34 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_35 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h23 == _T_1834) begin
          memory_35 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_36 <= 32'h8fc3001c;
    end else begin
      if (io_mem_wen) begin
        if (8'h24 == _T_1834) begin
          memory_36 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_37 <= 32'h24020008;
    end else begin
      if (io_mem_wen) begin
        if (8'h25 == _T_1834) begin
          memory_37 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_38 <= 32'h1462002e;
    end else begin
      if (io_mem_wen) begin
        if (8'h26 == _T_1834) begin
          memory_38 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_39 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h27 == _T_1834) begin
          memory_39 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_40 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h28 == _T_1834) begin
          memory_40 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_41 <= 32'h8c420350;
    end else begin
      if (io_mem_wen) begin
        if (8'h29 == _T_1834) begin
          memory_41 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_42 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h2a == _T_1834) begin
          memory_42 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_43 <= 32'h14400018;
    end else begin
      if (io_mem_wen) begin
        if (8'h2b == _T_1834) begin
          memory_43 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_44 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h2c == _T_1834) begin
          memory_44 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_45 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h2d == _T_1834) begin
          memory_45 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_46 <= 32'h24030018;
    end else begin
      if (io_mem_wen) begin
        if (8'h2e == _T_1834) begin
          memory_46 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_47 <= 32'hac430350;
    end else begin
      if (io_mem_wen) begin
        if (8'h2f == _T_1834) begin
          memory_47 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_48 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h30 == _T_1834) begin
          memory_48 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_49 <= 32'h8c420354;
    end else begin
      if (io_mem_wen) begin
        if (8'h31 == _T_1834) begin
          memory_49 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_50 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h32 == _T_1834) begin
          memory_50 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_51 <= 32'h2443ffff;
    end else begin
      if (io_mem_wen) begin
        if (8'h33 == _T_1834) begin
          memory_51 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_52 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h34 == _T_1834) begin
          memory_52 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_53 <= 32'hac430354;
    end else begin
      if (io_mem_wen) begin
        if (8'h35 == _T_1834) begin
          memory_53 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_54 <= 32'h24040f20;
    end else begin
      if (io_mem_wen) begin
        if (8'h36 == _T_1834) begin
          memory_54 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_55 <= 32'hc000076;
    end else begin
      if (io_mem_wen) begin
        if (8'h37 == _T_1834) begin
          memory_55 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_56 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h38 == _T_1834) begin
          memory_56 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_57 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h39 == _T_1834) begin
          memory_57 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_58 <= 32'h24030018;
    end else begin
      if (io_mem_wen) begin
        if (8'h3a == _T_1834) begin
          memory_58 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_59 <= 32'hac430350;
    end else begin
      if (io_mem_wen) begin
        if (8'h3b == _T_1834) begin
          memory_59 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_60 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h3c == _T_1834) begin
          memory_60 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_61 <= 32'h8c420354;
    end else begin
      if (io_mem_wen) begin
        if (8'h3d == _T_1834) begin
          memory_61 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_62 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h3e == _T_1834) begin
          memory_62 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_63 <= 32'h2443ffff;
    end else begin
      if (io_mem_wen) begin
        if (8'h3f == _T_1834) begin
          memory_63 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_64 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h40 == _T_1834) begin
          memory_64 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_65 <= 32'hac430354;
    end else begin
      if (io_mem_wen) begin
        if (8'h41 == _T_1834) begin
          memory_65 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_66 <= 32'h1000ffcc;
    end else begin
      if (io_mem_wen) begin
        if (8'h42 == _T_1834) begin
          memory_66 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_67 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h43 == _T_1834) begin
          memory_67 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_68 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h44 == _T_1834) begin
          memory_68 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_69 <= 32'h8c420350;
    end else begin
      if (io_mem_wen) begin
        if (8'h45 == _T_1834) begin
          memory_69 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_70 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h46 == _T_1834) begin
          memory_70 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_71 <= 32'h2443ffff;
    end else begin
      if (io_mem_wen) begin
        if (8'h47 == _T_1834) begin
          memory_71 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_72 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h48 == _T_1834) begin
          memory_72 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_73 <= 32'hac430350;
    end else begin
      if (io_mem_wen) begin
        if (8'h49 == _T_1834) begin
          memory_73 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_74 <= 32'h24040f20;
    end else begin
      if (io_mem_wen) begin
        if (8'h4a == _T_1834) begin
          memory_74 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_75 <= 32'hc000076;
    end else begin
      if (io_mem_wen) begin
        if (8'h4b == _T_1834) begin
          memory_75 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_76 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h4c == _T_1834) begin
          memory_76 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_77 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h4d == _T_1834) begin
          memory_77 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_78 <= 32'h8c420350;
    end else begin
      if (io_mem_wen) begin
        if (8'h4e == _T_1834) begin
          memory_78 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_79 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h4f == _T_1834) begin
          memory_79 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_80 <= 32'h2443ffff;
    end else begin
      if (io_mem_wen) begin
        if (8'h50 == _T_1834) begin
          memory_80 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_81 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h51 == _T_1834) begin
          memory_81 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_82 <= 32'hac430350;
    end else begin
      if (io_mem_wen) begin
        if (8'h52 == _T_1834) begin
          memory_82 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_83 <= 32'h1000ffbb;
    end else begin
      if (io_mem_wen) begin
        if (8'h53 == _T_1834) begin
          memory_83 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_84 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h54 == _T_1834) begin
          memory_84 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_85 <= 32'h8fc3001c;
    end else begin
      if (io_mem_wen) begin
        if (8'h55 == _T_1834) begin
          memory_85 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_86 <= 32'h2402001b;
    end else begin
      if (io_mem_wen) begin
        if (8'h56 == _T_1834) begin
          memory_86 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_87 <= 32'h14620016;
    end else begin
      if (io_mem_wen) begin
        if (8'h57 == _T_1834) begin
          memory_87 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_88 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h58 == _T_1834) begin
          memory_88 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_89 <= 32'hafc00018;
    end else begin
      if (io_mem_wen) begin
        if (8'h59 == _T_1834) begin
          memory_89 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_90 <= 32'h10000008;
    end else begin
      if (io_mem_wen) begin
        if (8'h5a == _T_1834) begin
          memory_90 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_91 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h5b == _T_1834) begin
          memory_91 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_92 <= 32'h24040f20;
    end else begin
      if (io_mem_wen) begin
        if (8'h5c == _T_1834) begin
          memory_92 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_93 <= 32'hc000076;
    end else begin
      if (io_mem_wen) begin
        if (8'h5d == _T_1834) begin
          memory_93 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_94 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h5e == _T_1834) begin
          memory_94 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_95 <= 32'h8fc20018;
    end else begin
      if (io_mem_wen) begin
        if (8'h5f == _T_1834) begin
          memory_95 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_96 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h60 == _T_1834) begin
          memory_96 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_97 <= 32'h24420001;
    end else begin
      if (io_mem_wen) begin
        if (8'h61 == _T_1834) begin
          memory_97 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_98 <= 32'hafc20018;
    end else begin
      if (io_mem_wen) begin
        if (8'h62 == _T_1834) begin
          memory_98 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_99 <= 32'h8fc20018;
    end else begin
      if (io_mem_wen) begin
        if (8'h63 == _T_1834) begin
          memory_99 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_100 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h64 == _T_1834) begin
          memory_100 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_101 <= 32'h28420fa0;
    end else begin
      if (io_mem_wen) begin
        if (8'h65 == _T_1834) begin
          memory_101 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_102 <= 32'h1440fff5;
    end else begin
      if (io_mem_wen) begin
        if (8'h66 == _T_1834) begin
          memory_102 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_103 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h67 == _T_1834) begin
          memory_103 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_104 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h68 == _T_1834) begin
          memory_104 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_105 <= 32'hac400350;
    end else begin
      if (io_mem_wen) begin
        if (8'h69 == _T_1834) begin
          memory_105 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_106 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h6a == _T_1834) begin
          memory_106 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_107 <= 32'hac400354;
    end else begin
      if (io_mem_wen) begin
        if (8'h6b == _T_1834) begin
          memory_107 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_108 <= 32'h1000ffa2;
    end else begin
      if (io_mem_wen) begin
        if (8'h6c == _T_1834) begin
          memory_108 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_109 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h6d == _T_1834) begin
          memory_109 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_110 <= 32'h8fc2001c;
    end else begin
      if (io_mem_wen) begin
        if (8'h6e == _T_1834) begin
          memory_110 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_111 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h6f == _T_1834) begin
          memory_111 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_112 <= 32'h34420f00;
    end else begin
      if (io_mem_wen) begin
        if (8'h70 == _T_1834) begin
          memory_112 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_113 <= 32'h402025;
    end else begin
      if (io_mem_wen) begin
        if (8'h71 == _T_1834) begin
          memory_113 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_114 <= 32'hc000076;
    end else begin
      if (io_mem_wen) begin
        if (8'h72 == _T_1834) begin
          memory_114 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_115 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h73 == _T_1834) begin
          memory_115 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_116 <= 32'h1000ff9a;
    end else begin
      if (io_mem_wen) begin
        if (8'h74 == _T_1834) begin
          memory_116 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_117 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h75 == _T_1834) begin
          memory_117 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_118 <= 32'h27bdffe8;
    end else begin
      if (io_mem_wen) begin
        if (8'h76 == _T_1834) begin
          memory_118 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_119 <= 32'hafbe0014;
    end else begin
      if (io_mem_wen) begin
        if (8'h77 == _T_1834) begin
          memory_119 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_120 <= 32'h3a0f025;
    end else begin
      if (io_mem_wen) begin
        if (8'h78 == _T_1834) begin
          memory_120 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_121 <= 32'hafc40018;
    end else begin
      if (io_mem_wen) begin
        if (8'h79 == _T_1834) begin
          memory_121 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_122 <= 32'h24023000;
    end else begin
      if (io_mem_wen) begin
        if (8'h7a == _T_1834) begin
          memory_122 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_123 <= 32'hafc20008;
    end else begin
      if (io_mem_wen) begin
        if (8'h7b == _T_1834) begin
          memory_123 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_124 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h7c == _T_1834) begin
          memory_124 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_125 <= 32'h8c430354;
    end else begin
      if (io_mem_wen) begin
        if (8'h7d == _T_1834) begin
          memory_125 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_126 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h7e == _T_1834) begin
          memory_126 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_127 <= 32'h601025;
    end else begin
      if (io_mem_wen) begin
        if (8'h7f == _T_1834) begin
          memory_127 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_128 <= 32'h21080;
    end else begin
      if (io_mem_wen) begin
        if (8'h80 == _T_1834) begin
          memory_128 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_129 <= 32'h431021;
    end else begin
      if (io_mem_wen) begin
        if (8'h81 == _T_1834) begin
          memory_129 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_130 <= 32'h21100;
    end else begin
      if (io_mem_wen) begin
        if (8'h82 == _T_1834) begin
          memory_130 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_131 <= 32'h401825;
    end else begin
      if (io_mem_wen) begin
        if (8'h83 == _T_1834) begin
          memory_131 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_132 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h84 == _T_1834) begin
          memory_132 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_133 <= 32'h8c420350;
    end else begin
      if (io_mem_wen) begin
        if (8'h85 == _T_1834) begin
          memory_133 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_134 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h86 == _T_1834) begin
          memory_134 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_135 <= 32'h621021;
    end else begin
      if (io_mem_wen) begin
        if (8'h87 == _T_1834) begin
          memory_135 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_136 <= 32'h21080;
    end else begin
      if (io_mem_wen) begin
        if (8'h88 == _T_1834) begin
          memory_136 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_137 <= 32'h8fc30008;
    end else begin
      if (io_mem_wen) begin
        if (8'h89 == _T_1834) begin
          memory_137 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_138 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h8a == _T_1834) begin
          memory_138 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_139 <= 32'h621021;
    end else begin
      if (io_mem_wen) begin
        if (8'h8b == _T_1834) begin
          memory_139 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_140 <= 32'h8fc30018;
    end else begin
      if (io_mem_wen) begin
        if (8'h8c == _T_1834) begin
          memory_140 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_141 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h8d == _T_1834) begin
          memory_141 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_142 <= 32'hac430000;
    end else begin
      if (io_mem_wen) begin
        if (8'h8e == _T_1834) begin
          memory_142 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_143 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h8f == _T_1834) begin
          memory_143 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_144 <= 32'h8c420350;
    end else begin
      if (io_mem_wen) begin
        if (8'h90 == _T_1834) begin
          memory_144 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_145 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h91 == _T_1834) begin
          memory_145 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_146 <= 32'h24430001;
    end else begin
      if (io_mem_wen) begin
        if (8'h92 == _T_1834) begin
          memory_146 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_147 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h93 == _T_1834) begin
          memory_147 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_148 <= 32'hac430350;
    end else begin
      if (io_mem_wen) begin
        if (8'h94 == _T_1834) begin
          memory_148 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_149 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h95 == _T_1834) begin
          memory_149 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_150 <= 32'h8c430350;
    end else begin
      if (io_mem_wen) begin
        if (8'h96 == _T_1834) begin
          memory_150 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_151 <= 32'h24020050;
    end else begin
      if (io_mem_wen) begin
        if (8'h97 == _T_1834) begin
          memory_151 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_152 <= 32'h14620010;
    end else begin
      if (io_mem_wen) begin
        if (8'h98 == _T_1834) begin
          memory_152 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_153 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h99 == _T_1834) begin
          memory_153 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_154 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h9a == _T_1834) begin
          memory_154 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_155 <= 32'hac400350;
    end else begin
      if (io_mem_wen) begin
        if (8'h9b == _T_1834) begin
          memory_155 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_156 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'h9c == _T_1834) begin
          memory_156 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_157 <= 32'h8c420354;
    end else begin
      if (io_mem_wen) begin
        if (8'h9d == _T_1834) begin
          memory_157 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_158 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'h9e == _T_1834) begin
          memory_158 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_159 <= 32'h24430001;
    end else begin
      if (io_mem_wen) begin
        if (8'h9f == _T_1834) begin
          memory_159 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_160 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'ha0 == _T_1834) begin
          memory_160 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_161 <= 32'hac430354;
    end else begin
      if (io_mem_wen) begin
        if (8'ha1 == _T_1834) begin
          memory_161 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_162 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'ha2 == _T_1834) begin
          memory_162 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_163 <= 32'h8c430354;
    end else begin
      if (io_mem_wen) begin
        if (8'ha3 == _T_1834) begin
          memory_163 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_164 <= 32'h24020019;
    end else begin
      if (io_mem_wen) begin
        if (8'ha4 == _T_1834) begin
          memory_164 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_165 <= 32'h14620003;
    end else begin
      if (io_mem_wen) begin
        if (8'ha5 == _T_1834) begin
          memory_165 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_166 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'ha6 == _T_1834) begin
          memory_166 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_167 <= 32'h3c020000;
    end else begin
      if (io_mem_wen) begin
        if (8'ha7 == _T_1834) begin
          memory_167 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_168 <= 32'hac400354;
    end else begin
      if (io_mem_wen) begin
        if (8'ha8 == _T_1834) begin
          memory_168 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_169 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'ha9 == _T_1834) begin
          memory_169 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_170 <= 32'h3c0e825;
    end else begin
      if (io_mem_wen) begin
        if (8'haa == _T_1834) begin
          memory_170 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_171 <= 32'h8fbe0014;
    end else begin
      if (io_mem_wen) begin
        if (8'hab == _T_1834) begin
          memory_171 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_172 <= 32'h27bd0018;
    end else begin
      if (io_mem_wen) begin
        if (8'hac == _T_1834) begin
          memory_172 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_173 <= 32'h3e00008;
    end else begin
      if (io_mem_wen) begin
        if (8'had == _T_1834) begin
          memory_173 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_174 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hae == _T_1834) begin
          memory_174 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_175 <= 32'h27bdffe0;
    end else begin
      if (io_mem_wen) begin
        if (8'haf == _T_1834) begin
          memory_175 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_176 <= 32'hafbe001c;
    end else begin
      if (io_mem_wen) begin
        if (8'hb0 == _T_1834) begin
          memory_176 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_177 <= 32'h3a0f025;
    end else begin
      if (io_mem_wen) begin
        if (8'hb1 == _T_1834) begin
          memory_177 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_178 <= 32'h3402ff00;
    end else begin
      if (io_mem_wen) begin
        if (8'hb2 == _T_1834) begin
          memory_178 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_179 <= 32'hafc20008;
    end else begin
      if (io_mem_wen) begin
        if (8'hb3 == _T_1834) begin
          memory_179 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_180 <= 32'h3c024000;
    end else begin
      if (io_mem_wen) begin
        if (8'hb4 == _T_1834) begin
          memory_180 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_181 <= 32'hafc2000c;
    end else begin
      if (io_mem_wen) begin
        if (8'hb5 == _T_1834) begin
          memory_181 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_182 <= 32'h240200ff;
    end else begin
      if (io_mem_wen) begin
        if (8'hb6 == _T_1834) begin
          memory_182 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_183 <= 32'hafc20010;
    end else begin
      if (io_mem_wen) begin
        if (8'hb7 == _T_1834) begin
          memory_183 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_184 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hb8 == _T_1834) begin
          memory_184 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_185 <= 32'h8fc20008;
    end else begin
      if (io_mem_wen) begin
        if (8'hb9 == _T_1834) begin
          memory_185 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_186 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hba == _T_1834) begin
          memory_186 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_187 <= 32'h8c430000;
    end else begin
      if (io_mem_wen) begin
        if (8'hbb == _T_1834) begin
          memory_187 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_188 <= 32'h8fc2000c;
    end else begin
      if (io_mem_wen) begin
        if (8'hbc == _T_1834) begin
          memory_188 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_189 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hbd == _T_1834) begin
          memory_189 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_190 <= 32'h621024;
    end else begin
      if (io_mem_wen) begin
        if (8'hbe == _T_1834) begin
          memory_190 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_191 <= 32'h1040fff9;
    end else begin
      if (io_mem_wen) begin
        if (8'hbf == _T_1834) begin
          memory_191 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_192 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hc0 == _T_1834) begin
          memory_192 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_193 <= 32'h8fc20008;
    end else begin
      if (io_mem_wen) begin
        if (8'hc1 == _T_1834) begin
          memory_193 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_194 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hc2 == _T_1834) begin
          memory_194 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_195 <= 32'h8c420000;
    end else begin
      if (io_mem_wen) begin
        if (8'hc3 == _T_1834) begin
          memory_195 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_196 <= 32'h8fc30010;
    end else begin
      if (io_mem_wen) begin
        if (8'hc4 == _T_1834) begin
          memory_196 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_197 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hc5 == _T_1834) begin
          memory_197 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_198 <= 32'h621024;
    end else begin
      if (io_mem_wen) begin
        if (8'hc6 == _T_1834) begin
          memory_198 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_199 <= 32'hafc20014;
    end else begin
      if (io_mem_wen) begin
        if (8'hc7 == _T_1834) begin
          memory_199 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_200 <= 32'h8fc20008;
    end else begin
      if (io_mem_wen) begin
        if (8'hc8 == _T_1834) begin
          memory_200 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_201 <= 32'h3c038000;
    end else begin
      if (io_mem_wen) begin
        if (8'hc9 == _T_1834) begin
          memory_201 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_202 <= 32'hac430000;
    end else begin
      if (io_mem_wen) begin
        if (8'hca == _T_1834) begin
          memory_202 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_203 <= 32'h8fc20014;
    end else begin
      if (io_mem_wen) begin
        if (8'hcb == _T_1834) begin
          memory_203 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_204 <= 32'h3c0e825;
    end else begin
      if (io_mem_wen) begin
        if (8'hcc == _T_1834) begin
          memory_204 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_205 <= 32'h8fbe001c;
    end else begin
      if (io_mem_wen) begin
        if (8'hcd == _T_1834) begin
          memory_205 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_206 <= 32'h27bd0020;
    end else begin
      if (io_mem_wen) begin
        if (8'hce == _T_1834) begin
          memory_206 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_207 <= 32'h3e00008;
    end else begin
      if (io_mem_wen) begin
        if (8'hcf == _T_1834) begin
          memory_207 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_208 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hd0 == _T_1834) begin
          memory_208 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_209 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hd1 == _T_1834) begin
          memory_209 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_210 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hd2 == _T_1834) begin
          memory_210 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_211 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hd3 == _T_1834) begin
          memory_211 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_212 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hd4 == _T_1834) begin
          memory_212 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_213 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hd5 == _T_1834) begin
          memory_213 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_214 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hd6 == _T_1834) begin
          memory_214 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_215 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hd7 == _T_1834) begin
          memory_215 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_216 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hd8 == _T_1834) begin
          memory_216 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_217 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hd9 == _T_1834) begin
          memory_217 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_218 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hda == _T_1834) begin
          memory_218 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_219 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hdb == _T_1834) begin
          memory_219 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_220 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hdc == _T_1834) begin
          memory_220 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_221 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hdd == _T_1834) begin
          memory_221 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_222 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hde == _T_1834) begin
          memory_222 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_223 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hdf == _T_1834) begin
          memory_223 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_224 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'he0 == _T_1834) begin
          memory_224 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_225 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'he1 == _T_1834) begin
          memory_225 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_226 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'he2 == _T_1834) begin
          memory_226 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_227 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'he3 == _T_1834) begin
          memory_227 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_228 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'he4 == _T_1834) begin
          memory_228 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_229 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'he5 == _T_1834) begin
          memory_229 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_230 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'he6 == _T_1834) begin
          memory_230 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_231 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'he7 == _T_1834) begin
          memory_231 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_232 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'he8 == _T_1834) begin
          memory_232 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_233 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'he9 == _T_1834) begin
          memory_233 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_234 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hea == _T_1834) begin
          memory_234 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_235 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'heb == _T_1834) begin
          memory_235 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_236 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hec == _T_1834) begin
          memory_236 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_237 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hed == _T_1834) begin
          memory_237 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_238 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hee == _T_1834) begin
          memory_238 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_239 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hef == _T_1834) begin
          memory_239 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_240 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hf0 == _T_1834) begin
          memory_240 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_241 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hf1 == _T_1834) begin
          memory_241 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_242 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hf2 == _T_1834) begin
          memory_242 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_243 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hf3 == _T_1834) begin
          memory_243 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_244 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hf4 == _T_1834) begin
          memory_244 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_245 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hf5 == _T_1834) begin
          memory_245 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_246 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hf6 == _T_1834) begin
          memory_246 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_247 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hf7 == _T_1834) begin
          memory_247 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_248 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hf8 == _T_1834) begin
          memory_248 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_249 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hf9 == _T_1834) begin
          memory_249 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_250 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hfa == _T_1834) begin
          memory_250 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_251 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hfb == _T_1834) begin
          memory_251 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_252 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hfc == _T_1834) begin
          memory_252 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_253 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hfd == _T_1834) begin
          memory_253 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_254 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hfe == _T_1834) begin
          memory_254 <= io_mem_wdata;
        end
      end
    end
    if (reset) begin
      memory_255 <= 32'h0;
    end else begin
      if (io_mem_wen) begin
        if (8'hff == _T_1834) begin
          memory_255 <= io_mem_wdata;
        end
      end
    end
  end
endmodule
module VGACore( // @[:@1122.2]
  input         clock, // @[:@1123.4]
  input         reset, // @[:@1124.4]
  output [31:0] io_row, // @[:@1125.4]
  output [31:0] io_col, // @[:@1125.4]
  output        io_ready, // @[:@1125.4]
  input  [11:0] io_color, // @[:@1125.4]
  output [3:0]  io_sig_r, // @[:@1125.4]
  output [3:0]  io_sig_g, // @[:@1125.4]
  output [3:0]  io_sig_b, // @[:@1125.4]
  output        io_sig_hsync, // @[:@1125.4]
  output        io_sig_vsync // @[:@1125.4]
);
  reg [31:0] h_tick; // @[VGACore.scala 136:23:@1127.4]
  reg [31:0] _RAND_0;
  reg [31:0] v_tick; // @[VGACore.scala 137:23:@1128.4]
  reg [31:0] _RAND_1;
  wire [32:0] _T_40; // @[VGACore.scala 143:25:@1141.4]
  wire [32:0] _T_41; // @[VGACore.scala 143:25:@1142.4]
  wire [31:0] _T_42; // @[VGACore.scala 143:25:@1143.4]
  wire  _T_43; // @[VGACore.scala 143:16:@1144.4]
  wire [32:0] _T_46; // @[VGACore.scala 145:27:@1147.6]
  wire [32:0] _T_47; // @[VGACore.scala 145:27:@1148.6]
  wire [31:0] _T_48; // @[VGACore.scala 145:27:@1149.6]
  wire  _T_49; // @[VGACore.scala 145:18:@1150.6]
  wire [32:0] _T_52; // @[VGACore.scala 148:24:@1155.8]
  wire [31:0] _T_53; // @[VGACore.scala 148:24:@1156.8]
  wire [31:0] _GEN_0; // @[VGACore.scala 145:34:@1151.6]
  wire [32:0] _T_55; // @[VGACore.scala 151:22:@1161.6]
  wire [31:0] _T_56; // @[VGACore.scala 151:22:@1162.6]
  wire [31:0] _GEN_1; // @[VGACore.scala 143:32:@1145.4]
  wire [31:0] _GEN_2; // @[VGACore.scala 143:32:@1145.4]
  wire  _T_59; // @[VGACore.scala 154:23:@1167.4]
  wire  _T_64; // @[VGACore.scala 154:46:@1172.4]
  wire  _T_65; // @[VGACore.scala 154:35:@1173.4]
  wire  _T_68; // @[VGACore.scala 154:73:@1176.4]
  wire  _T_69; // @[VGACore.scala 154:62:@1177.4]
  wire  _T_74; // @[VGACore.scala 154:96:@1182.4]
  wire [3:0] _T_111; // @[VGACore.scala 156:37:@1217.4]
  wire [3:0] _T_114; // @[VGACore.scala 157:37:@1220.4]
  wire [3:0] _T_117; // @[VGACore.scala 158:37:@1223.4]
  wire [32:0] _T_120; // @[VGACore.scala 160:20:@1226.4]
  wire [32:0] _T_121; // @[VGACore.scala 160:20:@1227.4]
  wire [31:0] _T_122; // @[VGACore.scala 160:20:@1228.4]
  wire [32:0] _T_123; // @[VGACore.scala 160:25:@1229.4]
  wire [32:0] _T_124; // @[VGACore.scala 160:25:@1230.4]
  wire [32:0] _T_126; // @[VGACore.scala 161:20:@1233.4]
  wire [32:0] _T_127; // @[VGACore.scala 161:20:@1234.4]
  wire [31:0] _T_128; // @[VGACore.scala 161:20:@1235.4]
  wire [32:0] _T_129; // @[VGACore.scala 161:25:@1236.4]
  wire [32:0] _T_130; // @[VGACore.scala 161:25:@1237.4]
  assign _T_40 = 32'h37e - 32'h1; // @[VGACore.scala 143:25:@1141.4]
  assign _T_41 = $unsigned(_T_40); // @[VGACore.scala 143:25:@1142.4]
  assign _T_42 = _T_41[31:0]; // @[VGACore.scala 143:25:@1143.4]
  assign _T_43 = h_tick >= _T_42; // @[VGACore.scala 143:16:@1144.4]
  assign _T_46 = 32'h1bd - 32'h1; // @[VGACore.scala 145:27:@1147.6]
  assign _T_47 = $unsigned(_T_46); // @[VGACore.scala 145:27:@1148.6]
  assign _T_48 = _T_47[31:0]; // @[VGACore.scala 145:27:@1149.6]
  assign _T_49 = v_tick >= _T_48; // @[VGACore.scala 145:18:@1150.6]
  assign _T_52 = v_tick + 32'h1; // @[VGACore.scala 148:24:@1155.8]
  assign _T_53 = v_tick + 32'h1; // @[VGACore.scala 148:24:@1156.8]
  assign _GEN_0 = _T_49 ? 32'h0 : _T_53; // @[VGACore.scala 145:34:@1151.6]
  assign _T_55 = h_tick + 32'h1; // @[VGACore.scala 151:22:@1161.6]
  assign _T_56 = h_tick + 32'h1; // @[VGACore.scala 151:22:@1162.6]
  assign _GEN_1 = _T_43 ? 32'h0 : _T_56; // @[VGACore.scala 143:32:@1145.4]
  assign _GEN_2 = _T_43 ? _GEN_0 : v_tick; // @[VGACore.scala 143:32:@1145.4]
  assign _T_59 = h_tick >= 32'h9f; // @[VGACore.scala 154:23:@1167.4]
  assign _T_64 = h_tick < 32'h36f; // @[VGACore.scala 154:46:@1172.4]
  assign _T_65 = _T_59 & _T_64; // @[VGACore.scala 154:35:@1173.4]
  assign _T_68 = v_tick >= 32'h22; // @[VGACore.scala 154:73:@1176.4]
  assign _T_69 = _T_65 & _T_68; // @[VGACore.scala 154:62:@1177.4]
  assign _T_74 = v_tick < 32'h1b2; // @[VGACore.scala 154:96:@1182.4]
  assign _T_111 = io_color[3:0]; // @[VGACore.scala 156:37:@1217.4]
  assign _T_114 = io_color[7:4]; // @[VGACore.scala 157:37:@1220.4]
  assign _T_117 = io_color[11:8]; // @[VGACore.scala 158:37:@1223.4]
  assign _T_120 = h_tick - 32'h6c; // @[VGACore.scala 160:20:@1226.4]
  assign _T_121 = $unsigned(_T_120); // @[VGACore.scala 160:20:@1227.4]
  assign _T_122 = _T_121[31:0]; // @[VGACore.scala 160:20:@1228.4]
  assign _T_123 = _T_122 - 32'h33; // @[VGACore.scala 160:25:@1229.4]
  assign _T_124 = $unsigned(_T_123); // @[VGACore.scala 160:25:@1230.4]
  assign _T_126 = v_tick - 32'h2; // @[VGACore.scala 161:20:@1233.4]
  assign _T_127 = $unsigned(_T_126); // @[VGACore.scala 161:20:@1234.4]
  assign _T_128 = _T_127[31:0]; // @[VGACore.scala 161:20:@1235.4]
  assign _T_129 = _T_128 - 32'h20; // @[VGACore.scala 161:25:@1236.4]
  assign _T_130 = $unsigned(_T_129); // @[VGACore.scala 161:25:@1237.4]
  assign io_row = _T_130[31:0]; // @[VGACore.scala 161:10:@1239.4]
  assign io_col = _T_124[31:0]; // @[VGACore.scala 160:10:@1232.4]
  assign io_ready = _T_69 & _T_74; // @[VGACore.scala 154:12:@1184.4]
  assign io_sig_r = io_ready ? _T_111 : 4'h0; // @[VGACore.scala 156:12:@1219.4]
  assign io_sig_g = io_ready ? _T_114 : 4'h0; // @[VGACore.scala 157:12:@1222.4]
  assign io_sig_b = io_ready ? _T_117 : 4'h0; // @[VGACore.scala 158:12:@1225.4]
  assign io_sig_hsync = h_tick >= 32'h6c; // @[VGACore.scala 163:16:@1241.4]
  assign io_sig_vsync = v_tick >= 32'h2; // @[VGACore.scala 164:16:@1243.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  h_tick = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  v_tick = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      h_tick <= 32'h0;
    end else begin
      if (_T_43) begin
        h_tick <= 32'h0;
      end else begin
        h_tick <= _T_56;
      end
    end
    if (reset) begin
      v_tick <= 32'h0;
    end else begin
      if (_T_43) begin
        if (_T_49) begin
          v_tick <= 32'h0;
        end else begin
          v_tick <= _T_53;
        end
      end
    end
  end
endmodule
module CGROM( // @[:@1254.2]
  input        clock, // @[:@1255.4]
  input  [7:0] io_addr, // @[:@1257.4]
  input  [3:0] io_row, // @[:@1257.4]
  output [7:0] io_data // @[:@1257.4]
);
  wire [7:0] impl_data; // @[VGA.scala 293:20:@1259.4]
  wire [3:0] impl_row; // @[VGA.scala 293:20:@1259.4]
  wire [7:0] impl_addr; // @[VGA.scala 293:20:@1259.4]
  wire  impl_clock; // @[VGA.scala 293:20:@1259.4]
  CGROMBlackbox impl ( // @[VGA.scala 293:20:@1259.4]
    .data(impl_data),
    .row(impl_row),
    .addr(impl_addr),
    .clock(impl_clock)
  );
  assign io_data = impl_data; // @[VGA.scala 297:11:@1267.4]
  assign impl_row = io_row; // @[VGA.scala 296:15:@1266.4]
  assign impl_addr = io_addr; // @[VGA.scala 295:16:@1265.4]
  assign impl_clock = clock; // @[VGA.scala 294:17:@1264.4]
endmodule
module VGA( // @[:@1269.2]
  input         clock, // @[:@1270.4]
  input         reset, // @[:@1271.4]
  output [3:0]  io_sig_r, // @[:@1272.4]
  output [3:0]  io_sig_g, // @[:@1272.4]
  output [3:0]  io_sig_b, // @[:@1272.4]
  output        io_sig_hsync, // @[:@1272.4]
  output        io_sig_vsync, // @[:@1272.4]
  output [31:0] io_vram_raddr, // @[:@1272.4]
  input  [15:0] io_vram_rdata // @[:@1272.4]
);
  wire  core_clock; // @[VGA.scala 156:20:@1274.4]
  wire  core_reset; // @[VGA.scala 156:20:@1274.4]
  wire [31:0] core_io_row; // @[VGA.scala 156:20:@1274.4]
  wire [31:0] core_io_col; // @[VGA.scala 156:20:@1274.4]
  wire  core_io_ready; // @[VGA.scala 156:20:@1274.4]
  wire [11:0] core_io_color; // @[VGA.scala 156:20:@1274.4]
  wire [3:0] core_io_sig_r; // @[VGA.scala 156:20:@1274.4]
  wire [3:0] core_io_sig_g; // @[VGA.scala 156:20:@1274.4]
  wire [3:0] core_io_sig_b; // @[VGA.scala 156:20:@1274.4]
  wire  core_io_sig_hsync; // @[VGA.scala 156:20:@1274.4]
  wire  core_io_sig_vsync; // @[VGA.scala 156:20:@1274.4]
  wire  cgrom_clock; // @[VGA.scala 157:21:@1277.4]
  wire [7:0] cgrom_io_addr; // @[VGA.scala 157:21:@1277.4]
  wire [3:0] cgrom_io_row; // @[VGA.scala 157:21:@1277.4]
  wire [7:0] cgrom_io_data; // @[VGA.scala 157:21:@1277.4]
  wire  _T_20; // @[VGA.scala 163:28:@1285.4]
  wire  _T_22; // @[VGA.scala 163:53:@1286.4]
  wire  start; // @[VGA.scala 163:37:@1287.4]
  reg [3:0] col_ctick; // @[Counter.scala 9:33:@1288.4]
  reg [31:0] _RAND_0;
  wire  _T_26; // @[Counter.scala 30:24:@1290.6]
  wire [4:0] _T_31; // @[Counter.scala 18:22:@1296.8]
  wire [3:0] _T_32; // @[Counter.scala 18:22:@1297.8]
  wire [3:0] _GEN_0; // @[Counter.scala 20:21:@1299.8]
  wire [3:0] _GEN_1; // @[Counter.scala 49:22:@1294.6]
  wire [3:0] _GEN_2; // @[Counter.scala 48:18:@1289.4]
  wire  col_ctick_carry; // @[Counter.scala 50:20:@1303.4]
  reg [6:0] col_tick; // @[Counter.scala 9:33:@1304.4]
  reg [31:0] _RAND_1;
  wire  _T_37; // @[Counter.scala 30:24:@1306.6]
  wire [7:0] _T_42; // @[Counter.scala 18:22:@1312.8]
  wire [6:0] _T_43; // @[Counter.scala 18:22:@1313.8]
  wire [6:0] _GEN_3; // @[Counter.scala 20:21:@1315.8]
  wire [6:0] _GEN_4; // @[Counter.scala 49:22:@1310.6]
  wire [6:0] _GEN_5; // @[Counter.scala 48:18:@1305.4]
  wire  col_tick_carry; // @[Counter.scala 50:20:@1319.4]
  reg [3:0] row_ctick; // @[Counter.scala 9:33:@1320.4]
  reg [31:0] _RAND_2;
  wire  _T_48; // @[Counter.scala 30:24:@1322.6]
  wire [4:0] _T_53; // @[Counter.scala 18:22:@1328.8]
  wire [3:0] _T_54; // @[Counter.scala 18:22:@1329.8]
  wire [3:0] _GEN_6; // @[Counter.scala 49:22:@1326.6]
  wire [3:0] _GEN_7; // @[Counter.scala 48:18:@1321.4]
  wire  row_ctick_carry; // @[Counter.scala 50:20:@1332.4]
  reg [4:0] row_tick; // @[Counter.scala 9:33:@1333.4]
  reg [31:0] _RAND_3;
  wire  _T_58; // @[Counter.scala 30:24:@1335.6]
  wire [5:0] _T_63; // @[Counter.scala 18:22:@1341.8]
  wire [4:0] _T_64; // @[Counter.scala 18:22:@1342.8]
  wire [4:0] _GEN_8; // @[Counter.scala 20:21:@1344.8]
  wire [4:0] _GEN_9; // @[Counter.scala 49:22:@1339.6]
  wire [4:0] _GEN_10; // @[Counter.scala 48:18:@1334.4]
  wire [2:0] _T_66; // @[VGA.scala 175:41:@1349.4]
  wire [3:0] _GEN_13; // @[Mux.scala 46:19:@1368.4]
  wire  _T_122; // @[Mux.scala 46:19:@1368.4]
  wire [11:0] _T_123; // @[Mux.scala 46:16:@1369.4]
  wire  _T_124; // @[Mux.scala 46:19:@1370.4]
  wire [11:0] _T_125; // @[Mux.scala 46:16:@1371.4]
  wire  _T_126; // @[Mux.scala 46:19:@1372.4]
  wire [11:0] _T_127; // @[Mux.scala 46:16:@1373.4]
  wire  _T_128; // @[Mux.scala 46:19:@1374.4]
  wire [11:0] _T_129; // @[Mux.scala 46:16:@1375.4]
  wire  _T_130; // @[Mux.scala 46:19:@1376.4]
  wire [11:0] _T_131; // @[Mux.scala 46:16:@1377.4]
  wire  _T_132; // @[Mux.scala 46:19:@1378.4]
  wire [11:0] _T_133; // @[Mux.scala 46:16:@1379.4]
  wire  _T_134; // @[Mux.scala 46:19:@1380.4]
  wire [11:0] _T_135; // @[Mux.scala 46:16:@1381.4]
  wire  _T_136; // @[Mux.scala 46:19:@1382.4]
  wire [11:0] _T_137; // @[Mux.scala 46:16:@1383.4]
  wire  _T_138; // @[Mux.scala 46:19:@1384.4]
  wire [11:0] bg_color; // @[Mux.scala 46:16:@1385.4]
  wire [3:0] _T_139; // @[VGA.scala 187:41:@1386.4]
  wire  _T_195; // @[Mux.scala 46:19:@1405.4]
  wire [11:0] _T_196; // @[Mux.scala 46:16:@1406.4]
  wire  _T_197; // @[Mux.scala 46:19:@1407.4]
  wire [11:0] _T_198; // @[Mux.scala 46:16:@1408.4]
  wire  _T_199; // @[Mux.scala 46:19:@1409.4]
  wire [11:0] _T_200; // @[Mux.scala 46:16:@1410.4]
  wire  _T_201; // @[Mux.scala 46:19:@1411.4]
  wire [11:0] _T_202; // @[Mux.scala 46:16:@1412.4]
  wire  _T_203; // @[Mux.scala 46:19:@1413.4]
  wire [11:0] _T_204; // @[Mux.scala 46:16:@1414.4]
  wire  _T_205; // @[Mux.scala 46:19:@1415.4]
  wire [11:0] _T_206; // @[Mux.scala 46:16:@1416.4]
  wire  _T_207; // @[Mux.scala 46:19:@1417.4]
  wire [11:0] _T_208; // @[Mux.scala 46:16:@1418.4]
  wire  _T_209; // @[Mux.scala 46:19:@1419.4]
  wire [11:0] _T_210; // @[Mux.scala 46:16:@1420.4]
  wire  _T_211; // @[Mux.scala 46:19:@1421.4]
  wire [11:0] fg_color; // @[Mux.scala 46:16:@1422.4]
  wire [31:0] _T_214; // @[VGA.scala 211:56:@1424.4]
  wire  _T_216; // @[VGA.scala 211:63:@1425.4]
  wire  frame_bp; // @[VGA.scala 211:40:@1426.4]
  wire [6:0] _GEN_14; // @[VGA.scala 212:33:@1427.4]
  wire [11:0] _T_218; // @[VGA.scala 212:33:@1427.4]
  wire [11:0] _GEN_15; // @[VGA.scala 212:40:@1428.4]
  wire [12:0] _T_219; // @[VGA.scala 212:40:@1428.4]
  wire [11:0] _T_220; // @[VGA.scala 212:40:@1429.4]
  wire [12:0] _T_222; // @[VGA.scala 212:51:@1430.4]
  wire [11:0] _T_223; // @[VGA.scala 212:51:@1431.4]
  wire  reach_the_end; // @[VGA.scala 212:57:@1432.4]
  wire [6:0] _GEN_18; // @[VGA.scala 218:46:@1443.8]
  wire [11:0] _T_237; // @[VGA.scala 218:46:@1443.8]
  wire  _T_239; // @[VGA.scala 218:53:@1444.8]
  wire [11:0] _T_246; // @[VGA.scala 218:28:@1448.8]
  wire [11:0] _GEN_11; // @[VGA.scala 217:31:@1440.6]
  wire [11:0] _T_257; // @[VGA.scala 223:26:@1462.6]
  wire [11:0] _GEN_12; // @[VGA.scala 216:28:@1438.4]
  wire  _T_259; // @[VGA.scala 226:35:@1465.4]
  wire  _T_261; // @[VGA.scala 226:46:@1466.4]
  wire  _T_262; // @[VGA.scala 226:43:@1467.4]
  wire  _T_264; // @[VGA.scala 228:17:@1468.4]
  wire  _T_267; // @[VGA.scala 229:6:@1469.4]
  wire [31:0] next_char_addr; // @[VGA.scala 215:28:@1436.4 VGA.scala 218:22:@1449.8 VGA.scala 220:22:@1453.8 VGA.scala 223:20:@1463.6]
  wire [31:0] _T_268; // @[Mux.scala 61:16:@1470.4]
  wire [31:0] _T_269; // @[Mux.scala 61:16:@1471.4]
  wire [7:0] _T_274; // @[VGA.scala 235:70:@1478.4]
  wire  _T_275; // @[VGA.scala 235:70:@1479.4]
  wire [11:0] _T_276; // @[VGA.scala 235:56:@1480.4]
  VGACore core ( // @[VGA.scala 156:20:@1274.4]
    .clock(core_clock),
    .reset(core_reset),
    .io_row(core_io_row),
    .io_col(core_io_col),
    .io_ready(core_io_ready),
    .io_color(core_io_color),
    .io_sig_r(core_io_sig_r),
    .io_sig_g(core_io_sig_g),
    .io_sig_b(core_io_sig_b),
    .io_sig_hsync(core_io_sig_hsync),
    .io_sig_vsync(core_io_sig_vsync)
  );
  CGROM cgrom ( // @[VGA.scala 157:21:@1277.4]
    .clock(cgrom_clock),
    .io_addr(cgrom_io_addr),
    .io_row(cgrom_io_row),
    .io_data(cgrom_io_data)
  );
  assign _T_20 = core_io_row == 32'h0; // @[VGA.scala 163:28:@1285.4]
  assign _T_22 = core_io_col == 32'h0; // @[VGA.scala 163:53:@1286.4]
  assign start = _T_20 & _T_22; // @[VGA.scala 163:37:@1287.4]
  assign _T_26 = col_ctick == 4'h8; // @[Counter.scala 30:24:@1290.6]
  assign _T_31 = col_ctick + 4'h1; // @[Counter.scala 18:22:@1296.8]
  assign _T_32 = col_ctick + 4'h1; // @[Counter.scala 18:22:@1297.8]
  assign _GEN_0 = _T_26 ? 4'h0 : _T_32; // @[Counter.scala 20:21:@1299.8]
  assign _GEN_1 = core_io_ready ? _GEN_0 : col_ctick; // @[Counter.scala 49:22:@1294.6]
  assign _GEN_2 = start ? 4'h1 : _GEN_1; // @[Counter.scala 48:18:@1289.4]
  assign col_ctick_carry = core_io_ready & _T_26; // @[Counter.scala 50:20:@1303.4]
  assign _T_37 = col_tick == 7'h4f; // @[Counter.scala 30:24:@1306.6]
  assign _T_42 = col_tick + 7'h1; // @[Counter.scala 18:22:@1312.8]
  assign _T_43 = col_tick + 7'h1; // @[Counter.scala 18:22:@1313.8]
  assign _GEN_3 = _T_37 ? 7'h0 : _T_43; // @[Counter.scala 20:21:@1315.8]
  assign _GEN_4 = col_ctick_carry ? _GEN_3 : col_tick; // @[Counter.scala 49:22:@1310.6]
  assign _GEN_5 = start ? 7'h0 : _GEN_4; // @[Counter.scala 48:18:@1305.4]
  assign col_tick_carry = col_ctick_carry & _T_37; // @[Counter.scala 50:20:@1319.4]
  assign _T_48 = row_ctick == 4'hf; // @[Counter.scala 30:24:@1322.6]
  assign _T_53 = row_ctick + 4'h1; // @[Counter.scala 18:22:@1328.8]
  assign _T_54 = row_ctick + 4'h1; // @[Counter.scala 18:22:@1329.8]
  assign _GEN_6 = col_tick_carry ? _T_54 : row_ctick; // @[Counter.scala 49:22:@1326.6]
  assign _GEN_7 = start ? 4'h0 : _GEN_6; // @[Counter.scala 48:18:@1321.4]
  assign row_ctick_carry = col_tick_carry & _T_48; // @[Counter.scala 50:20:@1332.4]
  assign _T_58 = row_tick == 5'h18; // @[Counter.scala 30:24:@1335.6]
  assign _T_63 = row_tick + 5'h1; // @[Counter.scala 18:22:@1341.8]
  assign _T_64 = row_tick + 5'h1; // @[Counter.scala 18:22:@1342.8]
  assign _GEN_8 = _T_58 ? 5'h0 : _T_64; // @[Counter.scala 20:21:@1344.8]
  assign _GEN_9 = row_ctick_carry ? _GEN_8 : row_tick; // @[Counter.scala 49:22:@1339.6]
  assign _GEN_10 = start ? 5'h0 : _GEN_9; // @[Counter.scala 48:18:@1334.4]
  assign _T_66 = io_vram_rdata[14:12]; // @[VGA.scala 175:41:@1349.4]
  assign _GEN_13 = {{1'd0}, _T_66}; // @[Mux.scala 46:19:@1368.4]
  assign _T_122 = 4'hf == _GEN_13; // @[Mux.scala 46:19:@1368.4]
  assign _T_123 = _T_122 ? 12'hfff : 12'h0; // @[Mux.scala 46:16:@1369.4]
  assign _T_124 = 3'h7 == _T_66; // @[Mux.scala 46:19:@1370.4]
  assign _T_125 = _T_124 ? 12'hccc : _T_123; // @[Mux.scala 46:16:@1371.4]
  assign _T_126 = 3'h6 == _T_66; // @[Mux.scala 46:19:@1372.4]
  assign _T_127 = _T_126 ? 12'hc60 : _T_125; // @[Mux.scala 46:16:@1373.4]
  assign _T_128 = 3'h5 == _T_66; // @[Mux.scala 46:19:@1374.4]
  assign _T_129 = _T_128 ? 12'hc0c : _T_127; // @[Mux.scala 46:16:@1375.4]
  assign _T_130 = 3'h4 == _T_66; // @[Mux.scala 46:19:@1376.4]
  assign _T_131 = _T_130 ? 12'hc00 : _T_129; // @[Mux.scala 46:16:@1377.4]
  assign _T_132 = 3'h3 == _T_66; // @[Mux.scala 46:19:@1378.4]
  assign _T_133 = _T_132 ? 12'hcc : _T_131; // @[Mux.scala 46:16:@1379.4]
  assign _T_134 = 3'h2 == _T_66; // @[Mux.scala 46:19:@1380.4]
  assign _T_135 = _T_134 ? 12'hc0 : _T_133; // @[Mux.scala 46:16:@1381.4]
  assign _T_136 = 3'h1 == _T_66; // @[Mux.scala 46:19:@1382.4]
  assign _T_137 = _T_136 ? 12'hc : _T_135; // @[Mux.scala 46:16:@1383.4]
  assign _T_138 = 3'h0 == _T_66; // @[Mux.scala 46:19:@1384.4]
  assign bg_color = _T_138 ? 12'h0 : _T_137; // @[Mux.scala 46:16:@1385.4]
  assign _T_139 = io_vram_rdata[11:8]; // @[VGA.scala 187:41:@1386.4]
  assign _T_195 = 4'hf == _T_139; // @[Mux.scala 46:19:@1405.4]
  assign _T_196 = _T_195 ? 12'hfff : 12'h0; // @[Mux.scala 46:16:@1406.4]
  assign _T_197 = 4'h7 == _T_139; // @[Mux.scala 46:19:@1407.4]
  assign _T_198 = _T_197 ? 12'hccc : _T_196; // @[Mux.scala 46:16:@1408.4]
  assign _T_199 = 4'h6 == _T_139; // @[Mux.scala 46:19:@1409.4]
  assign _T_200 = _T_199 ? 12'hc60 : _T_198; // @[Mux.scala 46:16:@1410.4]
  assign _T_201 = 4'h5 == _T_139; // @[Mux.scala 46:19:@1411.4]
  assign _T_202 = _T_201 ? 12'hc0c : _T_200; // @[Mux.scala 46:16:@1412.4]
  assign _T_203 = 4'h4 == _T_139; // @[Mux.scala 46:19:@1413.4]
  assign _T_204 = _T_203 ? 12'hc00 : _T_202; // @[Mux.scala 46:16:@1414.4]
  assign _T_205 = 4'h3 == _T_139; // @[Mux.scala 46:19:@1415.4]
  assign _T_206 = _T_205 ? 12'hcc : _T_204; // @[Mux.scala 46:16:@1416.4]
  assign _T_207 = 4'h2 == _T_139; // @[Mux.scala 46:19:@1417.4]
  assign _T_208 = _T_207 ? 12'hc0 : _T_206; // @[Mux.scala 46:16:@1418.4]
  assign _T_209 = 4'h1 == _T_139; // @[Mux.scala 46:19:@1419.4]
  assign _T_210 = _T_209 ? 12'hc : _T_208; // @[Mux.scala 46:16:@1420.4]
  assign _T_211 = 4'h0 == _T_139; // @[Mux.scala 46:19:@1421.4]
  assign fg_color = _T_211 ? 12'h0 : _T_210; // @[Mux.scala 46:16:@1422.4]
  assign _T_214 = $signed(core_io_col); // @[VGA.scala 211:56:@1424.4]
  assign _T_216 = $signed(_T_214) < $signed(32'sh0); // @[VGA.scala 211:63:@1425.4]
  assign frame_bp = _T_20 & _T_216; // @[VGA.scala 211:40:@1426.4]
  assign _GEN_14 = {{2'd0}, row_tick}; // @[VGA.scala 212:33:@1427.4]
  assign _T_218 = _GEN_14 * 7'h50; // @[VGA.scala 212:33:@1427.4]
  assign _GEN_15 = {{5'd0}, col_tick}; // @[VGA.scala 212:40:@1428.4]
  assign _T_219 = _T_218 + _GEN_15; // @[VGA.scala 212:40:@1428.4]
  assign _T_220 = _T_218 + _GEN_15; // @[VGA.scala 212:40:@1429.4]
  assign _T_222 = _T_220 + 12'h1; // @[VGA.scala 212:51:@1430.4]
  assign _T_223 = _T_220 + 12'h1; // @[VGA.scala 212:51:@1431.4]
  assign reach_the_end = _T_223 == 12'h7d0; // @[VGA.scala 212:57:@1432.4]
  assign _GEN_18 = {{2'd0}, _T_64}; // @[VGA.scala 218:46:@1443.8]
  assign _T_237 = _GEN_18 * 7'h50; // @[VGA.scala 218:46:@1443.8]
  assign _T_239 = _T_237 == 12'h7d0; // @[VGA.scala 218:53:@1444.8]
  assign _T_246 = _T_239 ? 12'h0 : _T_237; // @[VGA.scala 218:28:@1448.8]
  assign _GEN_11 = _T_48 ? _T_246 : _T_218; // @[VGA.scala 217:31:@1440.6]
  assign _T_257 = reach_the_end ? 12'h0 : _T_223; // @[VGA.scala 223:26:@1462.6]
  assign _GEN_12 = _T_37 ? _GEN_11 : _T_257; // @[VGA.scala 216:28:@1438.4]
  assign _T_259 = col_ctick != 4'h8; // @[VGA.scala 226:35:@1465.4]
  assign _T_261 = frame_bp == 1'h0; // @[VGA.scala 226:46:@1466.4]
  assign _T_262 = _T_259 & _T_261; // @[VGA.scala 226:43:@1467.4]
  assign _T_264 = frame_bp | reach_the_end; // @[VGA.scala 228:17:@1468.4]
  assign _T_267 = reach_the_end == 1'h0; // @[VGA.scala 229:6:@1469.4]
  assign next_char_addr = {{20'd0}, _GEN_12}; // @[VGA.scala 215:28:@1436.4 VGA.scala 218:22:@1449.8 VGA.scala 220:22:@1453.8 VGA.scala 223:20:@1463.6]
  assign _T_268 = _T_267 ? next_char_addr : 32'h0; // @[Mux.scala 61:16:@1470.4]
  assign _T_269 = _T_264 ? 32'h0 : _T_268; // @[Mux.scala 61:16:@1471.4]
  assign _T_274 = cgrom_io_data >> col_ctick; // @[VGA.scala 235:70:@1478.4]
  assign _T_275 = _T_274[0]; // @[VGA.scala 235:70:@1479.4]
  assign _T_276 = _T_275 ? fg_color : bg_color; // @[VGA.scala 235:56:@1480.4]
  assign io_sig_r = core_io_sig_r; // @[VGA.scala 159:15:@1284.4]
  assign io_sig_g = core_io_sig_g; // @[VGA.scala 159:15:@1283.4]
  assign io_sig_b = core_io_sig_b; // @[VGA.scala 159:15:@1282.4]
  assign io_sig_hsync = core_io_sig_hsync; // @[VGA.scala 159:15:@1281.4]
  assign io_sig_vsync = core_io_sig_vsync; // @[VGA.scala 159:15:@1280.4]
  assign io_vram_raddr = _T_262 ? {{20'd0}, _T_220} : _T_269; // @[VGA.scala 226:17:@1473.4]
  assign core_clock = clock; // @[:@1275.4]
  assign core_reset = reset; // @[:@1276.4]
  assign core_io_color = _T_26 ? bg_color : _T_276; // @[VGA.scala 235:17:@1482.4]
  assign cgrom_clock = clock; // @[:@1278.4]
  assign cgrom_io_addr = io_vram_rdata[7:0]; // @[VGA.scala 232:17:@1475.4]
  assign cgrom_io_row = row_ctick; // @[VGA.scala 233:17:@1476.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  col_ctick = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  col_tick = _RAND_1[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  row_ctick = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  row_tick = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      col_ctick <= 4'h0;
    end else begin
      if (start) begin
        col_ctick <= 4'h1;
      end else begin
        if (core_io_ready) begin
          if (_T_26) begin
            col_ctick <= 4'h0;
          end else begin
            col_ctick <= _T_32;
          end
        end
      end
    end
    if (reset) begin
      col_tick <= 7'h0;
    end else begin
      if (start) begin
        col_tick <= 7'h0;
      end else begin
        if (col_ctick_carry) begin
          if (_T_37) begin
            col_tick <= 7'h0;
          end else begin
            col_tick <= _T_43;
          end
        end
      end
    end
    if (reset) begin
      row_ctick <= 4'h0;
    end else begin
      if (start) begin
        row_ctick <= 4'h0;
      end else begin
        if (col_tick_carry) begin
          row_ctick <= _T_54;
        end
      end
    end
    if (reset) begin
      row_tick <= 5'h0;
    end else begin
      if (start) begin
        row_tick <= 5'h0;
      end else begin
        if (row_ctick_carry) begin
          if (_T_58) begin
            row_tick <= 5'h0;
          end else begin
            row_tick <= _T_64;
          end
        end
      end
    end
  end
endmodule
module DDU( // @[:@1484.2]
  input         clock, // @[:@1485.4]
  input         reset, // @[:@1486.4]
  input         io_cont, // @[:@1487.4]
  input         io_step, // @[:@1487.4]
  input         io_mem, // @[:@1487.4]
  input         io_inc, // @[:@1487.4]
  input         io_dec, // @[:@1487.4]
  output [6:0]  io_disp_seg, // @[:@1487.4]
  output        io_disp_dp, // @[:@1487.4]
  output [7:0]  io_disp_an, // @[:@1487.4]
  output [15:0] io_led, // @[:@1487.4]
  input  [15:0] io_vram_port_rdata, // @[:@1487.4]
  output [15:0] io_vram_port_raddr, // @[:@1487.4]
  output [15:0] io_vram_port_wdata, // @[:@1487.4]
  output [31:0] io_vram_port_waddr, // @[:@1487.4]
  output        io_vram_port_wen, // @[:@1487.4]
  input  [31:0] io_uart_port_mem_rdata, // @[:@1487.4]
  output [31:0] io_uart_port_mem_wdata, // @[:@1487.4]
  output        io_uart_port_mem_wen, // @[:@1487.4]
  output [3:0]  io_vga_sig_r, // @[:@1487.4]
  output [3:0]  io_vga_sig_g, // @[:@1487.4]
  output [3:0]  io_vga_sig_b, // @[:@1487.4]
  output        io_vga_sig_hsync, // @[:@1487.4]
  output        io_vga_sig_vsync // @[:@1487.4]
);
  wire  cpu_clock; // @[DDU.scala 41:21:@1489.4]
  wire  cpu_reset; // @[DDU.scala 41:21:@1489.4]
  wire [31:0] cpu_io_debug_pc; // @[DDU.scala 41:21:@1489.4]
  wire [4:0] cpu_io_debug_ra_c; // @[DDU.scala 41:21:@1489.4]
  wire [31:0] cpu_io_debug_rd_c; // @[DDU.scala 41:21:@1489.4]
  wire [31:0] cpu_io_debug_mr_a; // @[DDU.scala 41:21:@1489.4]
  wire [31:0] cpu_io_debug_mr_d; // @[DDU.scala 41:21:@1489.4]
  wire [31:0] cpu_io_mem_port_mem_rdata; // @[DDU.scala 41:21:@1489.4]
  wire [31:0] cpu_io_mem_port_mem_addr; // @[DDU.scala 41:21:@1489.4]
  wire [31:0] cpu_io_mem_port_mem_wdata; // @[DDU.scala 41:21:@1489.4]
  wire  cpu_io_mem_port_mem_wen; // @[DDU.scala 41:21:@1489.4]
  wire [31:0] cpu_io_mem_port_mem_addr2; // @[DDU.scala 41:21:@1489.4]
  wire [31:0] cpu_io_mem_port_mem_rdata2; // @[DDU.scala 41:21:@1489.4]
  wire  cpu_io_single; // @[DDU.scala 41:21:@1489.4]
  wire [31:0] mmap_io_mmap_port_mem_rdata; // @[DDU.scala 42:22:@1492.4]
  wire [31:0] mmap_io_mmap_port_mem_addr; // @[DDU.scala 42:22:@1492.4]
  wire [31:0] mmap_io_mmap_port_mem_wdata; // @[DDU.scala 42:22:@1492.4]
  wire  mmap_io_mmap_port_mem_wen; // @[DDU.scala 42:22:@1492.4]
  wire [31:0] mmap_io_mmap_port_mem_addr2; // @[DDU.scala 42:22:@1492.4]
  wire [31:0] mmap_io_mmap_port_mem_rdata2; // @[DDU.scala 42:22:@1492.4]
  wire [31:0] mmap_io_mem_port_mem_rdata; // @[DDU.scala 42:22:@1492.4]
  wire [31:0] mmap_io_mem_port_mem_addr; // @[DDU.scala 42:22:@1492.4]
  wire [31:0] mmap_io_mem_port_mem_wdata; // @[DDU.scala 42:22:@1492.4]
  wire  mmap_io_mem_port_mem_wen; // @[DDU.scala 42:22:@1492.4]
  wire [31:0] mmap_io_mem_port_mem_addr2; // @[DDU.scala 42:22:@1492.4]
  wire [31:0] mmap_io_mem_port_mem_rdata2; // @[DDU.scala 42:22:@1492.4]
  wire [31:0] mmap_io_uart_port_mem_rdata; // @[DDU.scala 42:22:@1492.4]
  wire [31:0] mmap_io_uart_port_mem_wdata; // @[DDU.scala 42:22:@1492.4]
  wire  mmap_io_uart_port_mem_wen; // @[DDU.scala 42:22:@1492.4]
  wire [31:0] mmap_io_vram_port_mem_addr; // @[DDU.scala 42:22:@1492.4]
  wire [15:0] mmap_io_vram_port_mem_wdata; // @[DDU.scala 42:22:@1492.4]
  wire  mmap_io_vram_port_mem_wen; // @[DDU.scala 42:22:@1492.4]
  wire  main_mem_clock; // @[DDU.scala 44:26:@1495.4]
  wire  main_mem_reset; // @[DDU.scala 44:26:@1495.4]
  wire [31:0] main_mem_io_mem_rdata; // @[DDU.scala 44:26:@1495.4]
  wire [31:0] main_mem_io_mem_addr; // @[DDU.scala 44:26:@1495.4]
  wire [31:0] main_mem_io_mem_wdata; // @[DDU.scala 44:26:@1495.4]
  wire  main_mem_io_mem_wen; // @[DDU.scala 44:26:@1495.4]
  wire [31:0] main_mem_io_mem_addr2; // @[DDU.scala 44:26:@1495.4]
  wire [31:0] main_mem_io_mem_rdata2; // @[DDU.scala 44:26:@1495.4]
  wire  vga_inst_clock; // @[DDU.scala 46:26:@1498.4]
  wire  vga_inst_reset; // @[DDU.scala 46:26:@1498.4]
  wire [3:0] vga_inst_io_sig_r; // @[DDU.scala 46:26:@1498.4]
  wire [3:0] vga_inst_io_sig_g; // @[DDU.scala 46:26:@1498.4]
  wire [3:0] vga_inst_io_sig_b; // @[DDU.scala 46:26:@1498.4]
  wire  vga_inst_io_sig_hsync; // @[DDU.scala 46:26:@1498.4]
  wire  vga_inst_io_sig_vsync; // @[DDU.scala 46:26:@1498.4]
  wire [31:0] vga_inst_io_vram_raddr; // @[DDU.scala 46:26:@1498.4]
  wire [15:0] vga_inst_io_vram_rdata; // @[DDU.scala 46:26:@1498.4]
  reg [12:0] _T_53; // @[DDU.scala 85:24:@1526.4]
  reg [31:0] _RAND_0;
  wire  _T_54; // @[DDU.scala 86:20:@1527.4]
  wire [13:0] _T_57; // @[DDU.scala 86:36:@1528.4]
  wire [12:0] _T_58; // @[DDU.scala 86:36:@1529.4]
  wire [12:0] _T_59; // @[DDU.scala 86:17:@1530.4]
  wire  _T_61; // @[DDU.scala 126:64:@1532.4]
  reg [2:0] step; // @[DDU.scala 91:24:@1533.4]
  reg [31:0] _RAND_1;
  wire  _T_64; // @[DDU.scala 92:31:@1534.4]
  wire [3:0] _T_67; // @[DDU.scala 92:47:@1535.4]
  wire [2:0] _T_68; // @[DDU.scala 92:47:@1536.4]
  wire [2:0] _T_69; // @[DDU.scala 92:28:@1537.4]
  wire [2:0] _T_70; // @[DDU.scala 92:17:@1538.4]
  wire [13:0] _T_72; // @[DDU.scala 127:30:@1540.4]
  wire [13:0] _T_73; // @[DDU.scala 127:19:@1541.4]
  wire [31:0] disp_data; // @[DDU.scala 144:21:@1602.4]
  wire [3:0] _T_77; // @[DDU.scala 132:25:@1544.4]
  wire [3:0] _T_79; // @[DDU.scala 133:25:@1545.4]
  wire [3:0] _T_81; // @[DDU.scala 134:25:@1546.4]
  wire [3:0] _T_83; // @[DDU.scala 135:25:@1547.4]
  wire [3:0] _T_85; // @[DDU.scala 136:25:@1548.4]
  wire [3:0] _T_87; // @[DDU.scala 137:25:@1549.4]
  wire [3:0] _T_89; // @[DDU.scala 138:25:@1550.4]
  wire [3:0] _T_91; // @[DDU.scala 139:25:@1551.4]
  wire  _T_92; // @[Mux.scala 46:19:@1552.4]
  wire [3:0] _T_93; // @[Mux.scala 46:16:@1553.4]
  wire  _T_94; // @[Mux.scala 46:19:@1554.4]
  wire [3:0] _T_95; // @[Mux.scala 46:16:@1555.4]
  wire  _T_96; // @[Mux.scala 46:19:@1556.4]
  wire [3:0] _T_97; // @[Mux.scala 46:16:@1557.4]
  wire  _T_98; // @[Mux.scala 46:19:@1558.4]
  wire [3:0] _T_99; // @[Mux.scala 46:16:@1559.4]
  wire  _T_100; // @[Mux.scala 46:19:@1560.4]
  wire [3:0] _T_101; // @[Mux.scala 46:16:@1561.4]
  wire  _T_102; // @[Mux.scala 46:19:@1562.4]
  wire [3:0] _T_103; // @[Mux.scala 46:16:@1563.4]
  wire  _T_104; // @[Mux.scala 46:19:@1564.4]
  wire [3:0] _T_105; // @[Mux.scala 46:16:@1565.4]
  wire  _T_106; // @[Mux.scala 46:19:@1566.4]
  wire [3:0] _T_107; // @[Mux.scala 46:16:@1567.4]
  wire  _T_141; // @[Mux.scala 46:19:@1568.4]
  wire [6:0] _T_142; // @[Mux.scala 46:16:@1569.4]
  wire  _T_143; // @[Mux.scala 46:19:@1570.4]
  wire [6:0] _T_144; // @[Mux.scala 46:16:@1571.4]
  wire  _T_145; // @[Mux.scala 46:19:@1572.4]
  wire [6:0] _T_146; // @[Mux.scala 46:16:@1573.4]
  wire  _T_147; // @[Mux.scala 46:19:@1574.4]
  wire [6:0] _T_148; // @[Mux.scala 46:16:@1575.4]
  wire  _T_149; // @[Mux.scala 46:19:@1576.4]
  wire [6:0] _T_150; // @[Mux.scala 46:16:@1577.4]
  wire  _T_151; // @[Mux.scala 46:19:@1578.4]
  wire [6:0] _T_152; // @[Mux.scala 46:16:@1579.4]
  wire  _T_153; // @[Mux.scala 46:19:@1580.4]
  wire [6:0] _T_154; // @[Mux.scala 46:16:@1581.4]
  wire  _T_155; // @[Mux.scala 46:19:@1582.4]
  wire [6:0] _T_156; // @[Mux.scala 46:16:@1583.4]
  wire  _T_157; // @[Mux.scala 46:19:@1584.4]
  wire [6:0] _T_158; // @[Mux.scala 46:16:@1585.4]
  wire  _T_159; // @[Mux.scala 46:19:@1586.4]
  wire [6:0] _T_160; // @[Mux.scala 46:16:@1587.4]
  wire  _T_161; // @[Mux.scala 46:19:@1588.4]
  wire [6:0] _T_162; // @[Mux.scala 46:16:@1589.4]
  wire  _T_163; // @[Mux.scala 46:19:@1590.4]
  wire [6:0] _T_164; // @[Mux.scala 46:16:@1591.4]
  wire  _T_165; // @[Mux.scala 46:19:@1592.4]
  wire [6:0] _T_166; // @[Mux.scala 46:16:@1593.4]
  wire  _T_167; // @[Mux.scala 46:19:@1594.4]
  wire [6:0] _T_168; // @[Mux.scala 46:16:@1595.4]
  wire  _T_169; // @[Mux.scala 46:19:@1596.4]
  wire [6:0] _T_170; // @[Mux.scala 46:16:@1597.4]
  wire  _T_171; // @[Mux.scala 46:19:@1598.4]
  reg [31:0] disp_addr; // @[DDU.scala 145:28:@1604.4]
  reg [31:0] _RAND_2;
  reg  _T_178; // @[DDU.scala 97:24:@1605.4]
  reg [31:0] _RAND_3;
  wire  _T_180; // @[DDU.scala 98:34:@1607.4]
  wire  _T_181; // @[DDU.scala 98:31:@1608.4]
  reg [21:0] _T_185; // @[DDU.scala 99:26:@1609.4]
  reg [31:0] _RAND_4;
  reg  _T_189; // @[DDU.scala 102:32:@1610.4]
  reg [31:0] _RAND_5;
  reg  _T_192; // @[DDU.scala 103:26:@1611.4]
  reg [31:0] _RAND_6;
  wire  _T_193; // @[DDU.scala 104:25:@1612.4]
  wire  _GEN_0; // @[DDU.scala 105:34:@1614.6]
  wire [21:0] _GEN_1; // @[DDU.scala 105:34:@1614.6]
  wire  _GEN_2; // @[DDU.scala 105:34:@1614.6]
  wire  _T_199; // @[DDU.scala 113:23:@1624.8]
  wire [22:0] _T_201; // @[DDU.scala 116:34:@1629.10]
  wire [22:0] _T_202; // @[DDU.scala 116:34:@1630.10]
  wire [21:0] _T_203; // @[DDU.scala 116:34:@1631.10]
  wire  _GEN_3; // @[DDU.scala 113:32:@1625.8]
  wire [21:0] _GEN_4; // @[DDU.scala 113:32:@1625.8]
  wire  _GEN_6; // @[DDU.scala 111:41:@1622.6]
  wire [21:0] _GEN_7; // @[DDU.scala 111:41:@1622.6]
  wire  _GEN_8; // @[DDU.scala 104:35:@1613.4]
  wire [21:0] _GEN_9; // @[DDU.scala 104:35:@1613.4]
  wire  _GEN_10; // @[DDU.scala 104:35:@1613.4]
  wire [32:0] _T_206; // @[DDU.scala 147:32:@1640.6]
  wire [31:0] _T_207; // @[DDU.scala 147:32:@1641.6]
  reg  _T_209; // @[DDU.scala 97:24:@1645.6]
  reg [31:0] _RAND_7;
  wire  _T_211; // @[DDU.scala 98:34:@1647.6]
  wire  _T_212; // @[DDU.scala 98:31:@1648.6]
  reg [21:0] _T_216; // @[DDU.scala 99:26:@1649.6]
  reg [31:0] _RAND_8;
  reg  _T_220; // @[DDU.scala 102:32:@1650.6]
  reg [31:0] _RAND_9;
  reg  _T_223; // @[DDU.scala 103:26:@1651.6]
  reg [31:0] _RAND_10;
  wire  _T_224; // @[DDU.scala 104:25:@1652.6]
  wire  _GEN_11; // @[DDU.scala 105:34:@1654.8]
  wire [21:0] _GEN_12; // @[DDU.scala 105:34:@1654.8]
  wire  _GEN_13; // @[DDU.scala 105:34:@1654.8]
  wire  _T_230; // @[DDU.scala 113:23:@1664.10]
  wire [22:0] _T_232; // @[DDU.scala 116:34:@1669.12]
  wire [22:0] _T_233; // @[DDU.scala 116:34:@1670.12]
  wire [21:0] _T_234; // @[DDU.scala 116:34:@1671.12]
  wire  _GEN_14; // @[DDU.scala 113:32:@1665.10]
  wire [21:0] _GEN_15; // @[DDU.scala 113:32:@1665.10]
  wire  _GEN_17; // @[DDU.scala 111:41:@1662.8]
  wire [21:0] _GEN_18; // @[DDU.scala 111:41:@1662.8]
  wire  _GEN_19; // @[DDU.scala 104:35:@1653.6]
  wire [21:0] _GEN_20; // @[DDU.scala 104:35:@1653.6]
  wire  _GEN_21; // @[DDU.scala 104:35:@1653.6]
  wire [32:0] _T_237; // @[DDU.scala 149:32:@1680.8]
  wire [32:0] _T_238; // @[DDU.scala 149:32:@1681.8]
  wire [31:0] _T_239; // @[DDU.scala 149:32:@1682.8]
  wire [31:0] _GEN_22; // @[DDU.scala 148:65:@1679.6]
  wire [31:0] _GEN_23; // @[DDU.scala 146:59:@1639.4]
  wire [4:0] _T_240; // @[DDU.scala 153:35:@1686.4]
  reg  _T_242; // @[DDU.scala 97:24:@1688.4]
  reg [31:0] _RAND_11;
  wire  _T_244; // @[DDU.scala 98:34:@1690.4]
  wire  _T_245; // @[DDU.scala 98:31:@1691.4]
  reg [21:0] _T_249; // @[DDU.scala 99:26:@1692.4]
  reg [31:0] _RAND_12;
  reg  _T_253; // @[DDU.scala 102:32:@1693.4]
  reg [31:0] _RAND_13;
  reg  pressed; // @[DDU.scala 103:26:@1694.4]
  reg [31:0] _RAND_14;
  wire  _T_256; // @[DDU.scala 104:25:@1695.4]
  wire  _GEN_24; // @[DDU.scala 105:34:@1697.6]
  wire [21:0] _GEN_25; // @[DDU.scala 105:34:@1697.6]
  wire  _GEN_26; // @[DDU.scala 105:34:@1697.6]
  wire  _T_262; // @[DDU.scala 113:23:@1707.8]
  wire [22:0] _T_264; // @[DDU.scala 116:34:@1712.10]
  wire [22:0] _T_265; // @[DDU.scala 116:34:@1713.10]
  wire [21:0] _T_266; // @[DDU.scala 116:34:@1714.10]
  wire  _GEN_27; // @[DDU.scala 113:32:@1708.8]
  wire [21:0] _GEN_28; // @[DDU.scala 113:32:@1708.8]
  wire  _GEN_30; // @[DDU.scala 111:41:@1705.6]
  wire [21:0] _GEN_31; // @[DDU.scala 111:41:@1705.6]
  wire  _GEN_32; // @[DDU.scala 104:35:@1696.4]
  wire [21:0] _GEN_33; // @[DDU.scala 104:35:@1696.4]
  wire  _GEN_34; // @[DDU.scala 104:35:@1696.4]
  wire  _T_268; // @[DDU.scala 158:32:@1722.4]
  wire [9:0] _T_271; // @[DDU.scala 164:42:@1725.4]
  wire [7:0] _T_272; // @[DDU.scala 164:48:@1726.4]
  wire [7:0] _T_274; // @[DDU.scala 164:24:@1728.4]
  wire [9:0] _T_275; // @[DDU.scala 164:89:@1729.4]
  wire [7:0] _T_276; // @[DDU.scala 164:95:@1730.4]
  CPU cpu ( // @[DDU.scala 41:21:@1489.4]
    .clock(cpu_clock),
    .reset(cpu_reset),
    .io_debug_pc(cpu_io_debug_pc),
    .io_debug_ra_c(cpu_io_debug_ra_c),
    .io_debug_rd_c(cpu_io_debug_rd_c),
    .io_debug_mr_a(cpu_io_debug_mr_a),
    .io_debug_mr_d(cpu_io_debug_mr_d),
    .io_mem_port_mem_rdata(cpu_io_mem_port_mem_rdata),
    .io_mem_port_mem_addr(cpu_io_mem_port_mem_addr),
    .io_mem_port_mem_wdata(cpu_io_mem_port_mem_wdata),
    .io_mem_port_mem_wen(cpu_io_mem_port_mem_wen),
    .io_mem_port_mem_addr2(cpu_io_mem_port_mem_addr2),
    .io_mem_port_mem_rdata2(cpu_io_mem_port_mem_rdata2),
    .io_single(cpu_io_single)
  );
  MMap mmap ( // @[DDU.scala 42:22:@1492.4]
    .io_mmap_port_mem_rdata(mmap_io_mmap_port_mem_rdata),
    .io_mmap_port_mem_addr(mmap_io_mmap_port_mem_addr),
    .io_mmap_port_mem_wdata(mmap_io_mmap_port_mem_wdata),
    .io_mmap_port_mem_wen(mmap_io_mmap_port_mem_wen),
    .io_mmap_port_mem_addr2(mmap_io_mmap_port_mem_addr2),
    .io_mmap_port_mem_rdata2(mmap_io_mmap_port_mem_rdata2),
    .io_mem_port_mem_rdata(mmap_io_mem_port_mem_rdata),
    .io_mem_port_mem_addr(mmap_io_mem_port_mem_addr),
    .io_mem_port_mem_wdata(mmap_io_mem_port_mem_wdata),
    .io_mem_port_mem_wen(mmap_io_mem_port_mem_wen),
    .io_mem_port_mem_addr2(mmap_io_mem_port_mem_addr2),
    .io_mem_port_mem_rdata2(mmap_io_mem_port_mem_rdata2),
    .io_uart_port_mem_rdata(mmap_io_uart_port_mem_rdata),
    .io_uart_port_mem_wdata(mmap_io_uart_port_mem_wdata),
    .io_uart_port_mem_wen(mmap_io_uart_port_mem_wen),
    .io_vram_port_mem_addr(mmap_io_vram_port_mem_addr),
    .io_vram_port_mem_wdata(mmap_io_vram_port_mem_wdata),
    .io_vram_port_mem_wen(mmap_io_vram_port_mem_wen)
  );
  Mem main_mem ( // @[DDU.scala 44:26:@1495.4]
    .clock(main_mem_clock),
    .reset(main_mem_reset),
    .io_mem_rdata(main_mem_io_mem_rdata),
    .io_mem_addr(main_mem_io_mem_addr),
    .io_mem_wdata(main_mem_io_mem_wdata),
    .io_mem_wen(main_mem_io_mem_wen),
    .io_mem_addr2(main_mem_io_mem_addr2),
    .io_mem_rdata2(main_mem_io_mem_rdata2)
  );
  VGA vga_inst ( // @[DDU.scala 46:26:@1498.4]
    .clock(vga_inst_clock),
    .reset(vga_inst_reset),
    .io_sig_r(vga_inst_io_sig_r),
    .io_sig_g(vga_inst_io_sig_g),
    .io_sig_b(vga_inst_io_sig_b),
    .io_sig_hsync(vga_inst_io_sig_hsync),
    .io_sig_vsync(vga_inst_io_sig_vsync),
    .io_vram_raddr(vga_inst_io_vram_raddr),
    .io_vram_rdata(vga_inst_io_vram_rdata)
  );
  assign _T_54 = _T_53 == 13'h1388; // @[DDU.scala 86:20:@1527.4]
  assign _T_57 = _T_53 + 13'h1; // @[DDU.scala 86:36:@1528.4]
  assign _T_58 = _T_53 + 13'h1; // @[DDU.scala 86:36:@1529.4]
  assign _T_59 = _T_54 ? 13'h0 : _T_58; // @[DDU.scala 86:17:@1530.4]
  assign _T_61 = _T_53 == 13'h0; // @[DDU.scala 126:64:@1532.4]
  assign _T_64 = step == 3'h7; // @[DDU.scala 92:31:@1534.4]
  assign _T_67 = step + 3'h1; // @[DDU.scala 92:47:@1535.4]
  assign _T_68 = step + 3'h1; // @[DDU.scala 92:47:@1536.4]
  assign _T_69 = _T_64 ? 3'h0 : _T_68; // @[DDU.scala 92:28:@1537.4]
  assign _T_70 = _T_61 ? _T_69 : step; // @[DDU.scala 92:17:@1538.4]
  assign _T_72 = 14'h1 << step; // @[DDU.scala 127:30:@1540.4]
  assign _T_73 = ~ _T_72; // @[DDU.scala 127:19:@1541.4]
  assign disp_data = io_mem ? cpu_io_debug_mr_d : cpu_io_debug_rd_c; // @[DDU.scala 144:21:@1602.4]
  assign _T_77 = disp_data[3:0]; // @[DDU.scala 132:25:@1544.4]
  assign _T_79 = disp_data[7:4]; // @[DDU.scala 133:25:@1545.4]
  assign _T_81 = disp_data[11:8]; // @[DDU.scala 134:25:@1546.4]
  assign _T_83 = disp_data[15:12]; // @[DDU.scala 135:25:@1547.4]
  assign _T_85 = disp_data[19:16]; // @[DDU.scala 136:25:@1548.4]
  assign _T_87 = disp_data[23:20]; // @[DDU.scala 137:25:@1549.4]
  assign _T_89 = disp_data[27:24]; // @[DDU.scala 138:25:@1550.4]
  assign _T_91 = disp_data[31:28]; // @[DDU.scala 139:25:@1551.4]
  assign _T_92 = 3'h7 == step; // @[Mux.scala 46:19:@1552.4]
  assign _T_93 = _T_92 ? _T_91 : 4'h0; // @[Mux.scala 46:16:@1553.4]
  assign _T_94 = 3'h6 == step; // @[Mux.scala 46:19:@1554.4]
  assign _T_95 = _T_94 ? _T_89 : _T_93; // @[Mux.scala 46:16:@1555.4]
  assign _T_96 = 3'h5 == step; // @[Mux.scala 46:19:@1556.4]
  assign _T_97 = _T_96 ? _T_87 : _T_95; // @[Mux.scala 46:16:@1557.4]
  assign _T_98 = 3'h4 == step; // @[Mux.scala 46:19:@1558.4]
  assign _T_99 = _T_98 ? _T_85 : _T_97; // @[Mux.scala 46:16:@1559.4]
  assign _T_100 = 3'h3 == step; // @[Mux.scala 46:19:@1560.4]
  assign _T_101 = _T_100 ? _T_83 : _T_99; // @[Mux.scala 46:16:@1561.4]
  assign _T_102 = 3'h2 == step; // @[Mux.scala 46:19:@1562.4]
  assign _T_103 = _T_102 ? _T_81 : _T_101; // @[Mux.scala 46:16:@1563.4]
  assign _T_104 = 3'h1 == step; // @[Mux.scala 46:19:@1564.4]
  assign _T_105 = _T_104 ? _T_79 : _T_103; // @[Mux.scala 46:16:@1565.4]
  assign _T_106 = 3'h0 == step; // @[Mux.scala 46:19:@1566.4]
  assign _T_107 = _T_106 ? _T_77 : _T_105; // @[Mux.scala 46:16:@1567.4]
  assign _T_141 = 4'hf == _T_107; // @[Mux.scala 46:19:@1568.4]
  assign _T_142 = _T_141 ? 7'he : 7'h40; // @[Mux.scala 46:16:@1569.4]
  assign _T_143 = 4'he == _T_107; // @[Mux.scala 46:19:@1570.4]
  assign _T_144 = _T_143 ? 7'h6 : _T_142; // @[Mux.scala 46:16:@1571.4]
  assign _T_145 = 4'hd == _T_107; // @[Mux.scala 46:19:@1572.4]
  assign _T_146 = _T_145 ? 7'h21 : _T_144; // @[Mux.scala 46:16:@1573.4]
  assign _T_147 = 4'hc == _T_107; // @[Mux.scala 46:19:@1574.4]
  assign _T_148 = _T_147 ? 7'h46 : _T_146; // @[Mux.scala 46:16:@1575.4]
  assign _T_149 = 4'hb == _T_107; // @[Mux.scala 46:19:@1576.4]
  assign _T_150 = _T_149 ? 7'h3 : _T_148; // @[Mux.scala 46:16:@1577.4]
  assign _T_151 = 4'ha == _T_107; // @[Mux.scala 46:19:@1578.4]
  assign _T_152 = _T_151 ? 7'h8 : _T_150; // @[Mux.scala 46:16:@1579.4]
  assign _T_153 = 4'h9 == _T_107; // @[Mux.scala 46:19:@1580.4]
  assign _T_154 = _T_153 ? 7'h10 : _T_152; // @[Mux.scala 46:16:@1581.4]
  assign _T_155 = 4'h8 == _T_107; // @[Mux.scala 46:19:@1582.4]
  assign _T_156 = _T_155 ? 7'h0 : _T_154; // @[Mux.scala 46:16:@1583.4]
  assign _T_157 = 4'h7 == _T_107; // @[Mux.scala 46:19:@1584.4]
  assign _T_158 = _T_157 ? 7'h78 : _T_156; // @[Mux.scala 46:16:@1585.4]
  assign _T_159 = 4'h6 == _T_107; // @[Mux.scala 46:19:@1586.4]
  assign _T_160 = _T_159 ? 7'h2 : _T_158; // @[Mux.scala 46:16:@1587.4]
  assign _T_161 = 4'h5 == _T_107; // @[Mux.scala 46:19:@1588.4]
  assign _T_162 = _T_161 ? 7'h12 : _T_160; // @[Mux.scala 46:16:@1589.4]
  assign _T_163 = 4'h4 == _T_107; // @[Mux.scala 46:19:@1590.4]
  assign _T_164 = _T_163 ? 7'h19 : _T_162; // @[Mux.scala 46:16:@1591.4]
  assign _T_165 = 4'h3 == _T_107; // @[Mux.scala 46:19:@1592.4]
  assign _T_166 = _T_165 ? 7'h30 : _T_164; // @[Mux.scala 46:16:@1593.4]
  assign _T_167 = 4'h2 == _T_107; // @[Mux.scala 46:19:@1594.4]
  assign _T_168 = _T_167 ? 7'h24 : _T_166; // @[Mux.scala 46:16:@1595.4]
  assign _T_169 = 4'h1 == _T_107; // @[Mux.scala 46:19:@1596.4]
  assign _T_170 = _T_169 ? 7'h79 : _T_168; // @[Mux.scala 46:16:@1597.4]
  assign _T_171 = 4'h0 == _T_107; // @[Mux.scala 46:19:@1598.4]
  assign _T_180 = _T_178 == 1'h0; // @[DDU.scala 98:34:@1607.4]
  assign _T_181 = io_inc & _T_180; // @[DDU.scala 98:31:@1608.4]
  assign _T_193 = _T_189 == 1'h0; // @[DDU.scala 104:25:@1612.4]
  assign _GEN_0 = _T_181 ? 1'h1 : _T_189; // @[DDU.scala 105:34:@1614.6]
  assign _GEN_1 = _T_181 ? 22'h2625a0 : _T_185; // @[DDU.scala 105:34:@1614.6]
  assign _GEN_2 = _T_181 ? 1'h1 : _T_192; // @[DDU.scala 105:34:@1614.6]
  assign _T_199 = _T_185 == 22'h0; // @[DDU.scala 113:23:@1624.8]
  assign _T_201 = _T_185 - 22'h1; // @[DDU.scala 116:34:@1629.10]
  assign _T_202 = $unsigned(_T_201); // @[DDU.scala 116:34:@1630.10]
  assign _T_203 = _T_202[21:0]; // @[DDU.scala 116:34:@1631.10]
  assign _GEN_3 = _T_199 ? 1'h0 : _T_189; // @[DDU.scala 113:32:@1625.8]
  assign _GEN_4 = _T_199 ? _T_185 : _T_203; // @[DDU.scala 113:32:@1625.8]
  assign _GEN_6 = _T_189 ? _GEN_3 : 1'h0; // @[DDU.scala 111:41:@1622.6]
  assign _GEN_7 = _T_189 ? _GEN_4 : _T_185; // @[DDU.scala 111:41:@1622.6]
  assign _GEN_8 = _T_193 ? _GEN_0 : _GEN_6; // @[DDU.scala 104:35:@1613.4]
  assign _GEN_9 = _T_193 ? _GEN_1 : _GEN_7; // @[DDU.scala 104:35:@1613.4]
  assign _GEN_10 = _T_193 ? _GEN_2 : 1'h0; // @[DDU.scala 104:35:@1613.4]
  assign _T_206 = disp_addr + 32'h1; // @[DDU.scala 147:32:@1640.6]
  assign _T_207 = disp_addr + 32'h1; // @[DDU.scala 147:32:@1641.6]
  assign _T_211 = _T_209 == 1'h0; // @[DDU.scala 98:34:@1647.6]
  assign _T_212 = io_dec & _T_211; // @[DDU.scala 98:31:@1648.6]
  assign _T_224 = _T_220 == 1'h0; // @[DDU.scala 104:25:@1652.6]
  assign _GEN_11 = _T_212 ? 1'h1 : _T_220; // @[DDU.scala 105:34:@1654.8]
  assign _GEN_12 = _T_212 ? 22'h2625a0 : _T_216; // @[DDU.scala 105:34:@1654.8]
  assign _GEN_13 = _T_212 ? 1'h1 : _T_223; // @[DDU.scala 105:34:@1654.8]
  assign _T_230 = _T_216 == 22'h0; // @[DDU.scala 113:23:@1664.10]
  assign _T_232 = _T_216 - 22'h1; // @[DDU.scala 116:34:@1669.12]
  assign _T_233 = $unsigned(_T_232); // @[DDU.scala 116:34:@1670.12]
  assign _T_234 = _T_233[21:0]; // @[DDU.scala 116:34:@1671.12]
  assign _GEN_14 = _T_230 ? 1'h0 : _T_220; // @[DDU.scala 113:32:@1665.10]
  assign _GEN_15 = _T_230 ? _T_216 : _T_234; // @[DDU.scala 113:32:@1665.10]
  assign _GEN_17 = _T_220 ? _GEN_14 : 1'h0; // @[DDU.scala 111:41:@1662.8]
  assign _GEN_18 = _T_220 ? _GEN_15 : _T_216; // @[DDU.scala 111:41:@1662.8]
  assign _GEN_19 = _T_224 ? _GEN_11 : _GEN_17; // @[DDU.scala 104:35:@1653.6]
  assign _GEN_20 = _T_224 ? _GEN_12 : _GEN_18; // @[DDU.scala 104:35:@1653.6]
  assign _GEN_21 = _T_224 ? _GEN_13 : 1'h0; // @[DDU.scala 104:35:@1653.6]
  assign _T_237 = disp_addr - 32'h1; // @[DDU.scala 149:32:@1680.8]
  assign _T_238 = $unsigned(_T_237); // @[DDU.scala 149:32:@1681.8]
  assign _T_239 = _T_238[31:0]; // @[DDU.scala 149:32:@1682.8]
  assign _GEN_22 = _T_223 ? _T_239 : disp_addr; // @[DDU.scala 148:65:@1679.6]
  assign _GEN_23 = _T_192 ? _T_207 : _GEN_22; // @[DDU.scala 146:59:@1639.4]
  assign _T_240 = disp_addr[4:0]; // @[DDU.scala 153:35:@1686.4]
  assign _T_244 = _T_242 == 1'h0; // @[DDU.scala 98:34:@1690.4]
  assign _T_245 = io_step & _T_244; // @[DDU.scala 98:31:@1691.4]
  assign _T_256 = _T_253 == 1'h0; // @[DDU.scala 104:25:@1695.4]
  assign _GEN_24 = _T_245 ? 1'h1 : _T_253; // @[DDU.scala 105:34:@1697.6]
  assign _GEN_25 = _T_245 ? 22'h2625a0 : _T_249; // @[DDU.scala 105:34:@1697.6]
  assign _GEN_26 = _T_245 ? 1'h1 : pressed; // @[DDU.scala 105:34:@1697.6]
  assign _T_262 = _T_249 == 22'h0; // @[DDU.scala 113:23:@1707.8]
  assign _T_264 = _T_249 - 22'h1; // @[DDU.scala 116:34:@1712.10]
  assign _T_265 = $unsigned(_T_264); // @[DDU.scala 116:34:@1713.10]
  assign _T_266 = _T_265[21:0]; // @[DDU.scala 116:34:@1714.10]
  assign _GEN_27 = _T_262 ? 1'h0 : _T_253; // @[DDU.scala 113:32:@1708.8]
  assign _GEN_28 = _T_262 ? _T_249 : _T_266; // @[DDU.scala 113:32:@1708.8]
  assign _GEN_30 = _T_253 ? _GEN_27 : 1'h0; // @[DDU.scala 111:41:@1705.6]
  assign _GEN_31 = _T_253 ? _GEN_28 : _T_249; // @[DDU.scala 111:41:@1705.6]
  assign _GEN_32 = _T_256 ? _GEN_24 : _GEN_30; // @[DDU.scala 104:35:@1696.4]
  assign _GEN_33 = _T_256 ? _GEN_25 : _GEN_31; // @[DDU.scala 104:35:@1696.4]
  assign _GEN_34 = _T_256 ? _GEN_26 : 1'h0; // @[DDU.scala 104:35:@1696.4]
  assign _T_268 = pressed | io_cont; // @[DDU.scala 158:32:@1722.4]
  assign _T_271 = disp_addr[9:0]; // @[DDU.scala 164:42:@1725.4]
  assign _T_272 = _T_271[9:2]; // @[DDU.scala 164:48:@1726.4]
  assign _T_274 = io_mem ? _T_272 : {{3'd0}, _T_240}; // @[DDU.scala 164:24:@1728.4]
  assign _T_275 = cpu_io_debug_pc[9:0]; // @[DDU.scala 164:89:@1729.4]
  assign _T_276 = _T_275[9:2]; // @[DDU.scala 164:95:@1730.4]
  assign io_disp_seg = _T_171 ? 7'h40 : _T_170; // @[DDU.scala 131:17:@1600.4]
  assign io_disp_dp = 1'h0; // @[DDU.scala 142:16:@1601.4]
  assign io_disp_an = _T_73[7:0]; // @[DDU.scala 127:16:@1542.4]
  assign io_led = {_T_274,_T_276}; // @[DDU.scala 164:12:@1733.4]
  assign io_vram_port_raddr = vga_inst_io_vram_raddr[15:0]; // @[DDU.scala 55:24:@1522.4]
  assign io_vram_port_wdata = mmap_io_vram_port_mem_wdata; // @[DDU.scala 57:24:@1523.4]
  assign io_vram_port_waddr = mmap_io_vram_port_mem_addr; // @[DDU.scala 58:24:@1524.4]
  assign io_vram_port_wen = mmap_io_vram_port_mem_wen; // @[DDU.scala 59:24:@1525.4]
  assign io_uart_port_mem_wdata = mmap_io_uart_port_mem_wdata; // @[DDU.scala 50:23:@1514.4]
  assign io_uart_port_mem_wen = mmap_io_uart_port_mem_wen; // @[DDU.scala 50:23:@1513.4]
  assign io_vga_sig_r = vga_inst_io_sig_r; // @[DDU.scala 52:21:@1520.4]
  assign io_vga_sig_g = vga_inst_io_sig_g; // @[DDU.scala 52:21:@1519.4]
  assign io_vga_sig_b = vga_inst_io_sig_b; // @[DDU.scala 52:21:@1518.4]
  assign io_vga_sig_hsync = vga_inst_io_sig_hsync; // @[DDU.scala 52:21:@1517.4]
  assign io_vga_sig_vsync = vga_inst_io_sig_vsync; // @[DDU.scala 52:21:@1516.4]
  assign cpu_clock = clock; // @[:@1490.4]
  assign cpu_reset = reset; // @[:@1491.4]
  assign cpu_io_debug_ra_c = disp_addr[4:0]; // @[DDU.scala 153:23:@1687.4]
  assign cpu_io_debug_mr_a = disp_addr; // @[DDU.scala 152:23:@1685.4]
  assign cpu_io_mem_port_mem_rdata = mmap_io_mmap_port_mem_rdata; // @[DDU.scala 48:21:@1506.4]
  assign cpu_io_mem_port_mem_rdata2 = mmap_io_mmap_port_mem_rdata2; // @[DDU.scala 48:21:@1501.4]
  assign cpu_io_single = _T_268 == 1'h0; // @[DDU.scala 158:19:@1724.4]
  assign mmap_io_mmap_port_mem_addr = cpu_io_mem_port_mem_addr; // @[DDU.scala 48:21:@1505.4]
  assign mmap_io_mmap_port_mem_wdata = cpu_io_mem_port_mem_wdata; // @[DDU.scala 48:21:@1504.4]
  assign mmap_io_mmap_port_mem_wen = cpu_io_mem_port_mem_wen; // @[DDU.scala 48:21:@1503.4]
  assign mmap_io_mmap_port_mem_addr2 = cpu_io_mem_port_mem_addr2; // @[DDU.scala 48:21:@1502.4]
  assign mmap_io_mem_port_mem_rdata = main_mem_io_mem_rdata; // @[DDU.scala 49:22:@1512.4]
  assign mmap_io_mem_port_mem_rdata2 = main_mem_io_mem_rdata2; // @[DDU.scala 49:22:@1507.4]
  assign mmap_io_uart_port_mem_rdata = io_uart_port_mem_rdata; // @[DDU.scala 50:23:@1515.4]
  assign main_mem_clock = clock; // @[:@1496.4]
  assign main_mem_reset = reset; // @[:@1497.4]
  assign main_mem_io_mem_addr = mmap_io_mem_port_mem_addr; // @[DDU.scala 49:22:@1511.4]
  assign main_mem_io_mem_wdata = mmap_io_mem_port_mem_wdata; // @[DDU.scala 49:22:@1510.4]
  assign main_mem_io_mem_wen = mmap_io_mem_port_mem_wen; // @[DDU.scala 49:22:@1509.4]
  assign main_mem_io_mem_addr2 = mmap_io_mem_port_mem_addr2; // @[DDU.scala 49:22:@1508.4]
  assign vga_inst_clock = clock; // @[:@1499.4]
  assign vga_inst_reset = reset; // @[:@1500.4]
  assign vga_inst_io_vram_rdata = io_vram_port_rdata; // @[DDU.scala 54:29:@1521.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_53 = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  step = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  disp_addr = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_178 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_185 = _RAND_4[21:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_189 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_192 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_209 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_216 = _RAND_8[21:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_220 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_223 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_242 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_249 = _RAND_12[21:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_253 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  pressed = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_53 <= 13'h0;
    end else begin
      if (_T_54) begin
        _T_53 <= 13'h0;
      end else begin
        _T_53 <= _T_58;
      end
    end
    if (reset) begin
      step <= 3'h0;
    end else begin
      if (_T_61) begin
        if (_T_64) begin
          step <= 3'h0;
        end else begin
          step <= _T_68;
        end
      end
    end
    if (reset) begin
      disp_addr <= 32'h0;
    end else begin
      if (_T_192) begin
        disp_addr <= _T_207;
      end else begin
        if (_T_223) begin
          disp_addr <= _T_239;
        end
      end
    end
    _T_178 <= io_inc;
    if (reset) begin
      _T_185 <= 22'h0;
    end else begin
      if (_T_193) begin
        if (_T_181) begin
          _T_185 <= 22'h2625a0;
        end
      end else begin
        if (_T_189) begin
          if (!(_T_199)) begin
            _T_185 <= _T_203;
          end
        end
      end
    end
    if (reset) begin
      _T_189 <= 1'h0;
    end else begin
      if (_T_193) begin
        if (_T_181) begin
          _T_189 <= 1'h1;
        end
      end else begin
        if (_T_189) begin
          if (_T_199) begin
            _T_189 <= 1'h0;
          end
        end else begin
          _T_189 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_192 <= 1'h0;
    end else begin
      if (_T_193) begin
        if (_T_181) begin
          _T_192 <= 1'h1;
        end
      end else begin
        _T_192 <= 1'h0;
      end
    end
    _T_209 <= io_dec;
    if (reset) begin
      _T_216 <= 22'h0;
    end else begin
      if (_T_224) begin
        if (_T_212) begin
          _T_216 <= 22'h2625a0;
        end
      end else begin
        if (_T_220) begin
          if (!(_T_230)) begin
            _T_216 <= _T_234;
          end
        end
      end
    end
    if (reset) begin
      _T_220 <= 1'h0;
    end else begin
      if (_T_224) begin
        if (_T_212) begin
          _T_220 <= 1'h1;
        end
      end else begin
        if (_T_220) begin
          if (_T_230) begin
            _T_220 <= 1'h0;
          end
        end else begin
          _T_220 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_223 <= 1'h0;
    end else begin
      if (_T_224) begin
        if (_T_212) begin
          _T_223 <= 1'h1;
        end
      end else begin
        _T_223 <= 1'h0;
      end
    end
    _T_242 <= io_step;
    if (reset) begin
      _T_249 <= 22'h0;
    end else begin
      if (_T_256) begin
        if (_T_245) begin
          _T_249 <= 22'h2625a0;
        end
      end else begin
        if (_T_253) begin
          if (!(_T_262)) begin
            _T_249 <= _T_266;
          end
        end
      end
    end
    if (reset) begin
      _T_253 <= 1'h0;
    end else begin
      if (_T_256) begin
        if (_T_245) begin
          _T_253 <= 1'h1;
        end
      end else begin
        if (_T_253) begin
          if (_T_262) begin
            _T_253 <= 1'h0;
          end
        end else begin
          _T_253 <= 1'h0;
        end
      end
    end
    if (reset) begin
      pressed <= 1'h0;
    end else begin
      if (_T_256) begin
        if (_T_245) begin
          pressed <= 1'h1;
        end
      end else begin
        pressed <= 1'h0;
      end
    end
  end
endmodule
